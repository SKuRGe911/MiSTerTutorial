//VERILOG ROM

module
data_io_rom
(
	input		wire	[31:0]	address,
	input		wire				clock,
	output	reg	[15:0]	q=16'd0
);

always @(posedge clock) begin
	case(address)
		32'h00000000: begin
				q			<=			16'h400B;
		end
		32'h00000002: begin
				q			<=			16'h0800;
		end
		32'h00000004: begin
				q			<=			16'h600B;
		end
		32'h00000006: begin
				q			<=			16'h0600;
		end
		32'h00000008: begin
				q			<=			16'h006F;
		end
		32'h0000000A: begin
				q			<=			16'h3D80;
		end
		32'h0000000C: begin
				q			<=			16'h0013;
		end
		32'h0000000E: begin
				q			<=			16'h0000;
		end
		32'h00000010: begin
				q			<=			16'hA10B;
		end
		32'h00000012: begin
				q			<=			16'h0200;
		end
		32'h00000014: begin
				q			<=			16'h218B;
		end
		32'h00000016: begin
				q			<=			16'h0201;
		end
		32'h00000018: begin
				q			<=			16'h00B7;
		end
		32'h0000001A: begin
				q			<=			16'h0000;
		end
		32'h0000001C: begin
				q			<=			16'h8093;
		end
		32'h0000001E: begin
				q			<=			16'h1600;
		end
		32'h00000020: begin
				q			<=			16'h410B;
		end
		32'h00000022: begin
				q			<=			16'h0000;
		end
		32'h00000024: begin
				q			<=			16'hA023;
		end
		32'h00000026: begin
				q			<=			16'h0020;
		end
		32'h00000028: begin
				q			<=			16'h410B;
		end
		32'h0000002A: begin
				q			<=			16'h0001;
		end
		32'h0000002C: begin
				q			<=			16'hA223;
		end
		32'h0000002E: begin
				q			<=			16'h0020;
		end
		32'h00000030: begin
				q			<=			16'hC10B;
		end
		32'h00000032: begin
				q			<=			16'h0001;
		end
		32'h00000034: begin
				q			<=			16'hA423;
		end
		32'h00000036: begin
				q			<=			16'h0020;
		end
		32'h00000038: begin
				q			<=			16'hA623;
		end
		32'h0000003A: begin
				q			<=			16'h0030;
		end
		32'h0000003C: begin
				q			<=			16'hA823;
		end
		32'h0000003E: begin
				q			<=			16'h0040;
		end
		32'h00000040: begin
				q			<=			16'hAA23;
		end
		32'h00000042: begin
				q			<=			16'h0050;
		end
		32'h00000044: begin
				q			<=			16'hAC23;
		end
		32'h00000046: begin
				q			<=			16'h0060;
		end
		32'h00000048: begin
				q			<=			16'hAE23;
		end
		32'h0000004A: begin
				q			<=			16'h0070;
		end
		32'h0000004C: begin
				q			<=			16'hA023;
		end
		32'h0000004E: begin
				q			<=			16'h0280;
		end
		32'h00000050: begin
				q			<=			16'hA223;
		end
		32'h00000052: begin
				q			<=			16'h0290;
		end
		32'h00000054: begin
				q			<=			16'hA423;
		end
		32'h00000056: begin
				q			<=			16'h02A0;
		end
		32'h00000058: begin
				q			<=			16'hA623;
		end
		32'h0000005A: begin
				q			<=			16'h02B0;
		end
		32'h0000005C: begin
				q			<=			16'hA823;
		end
		32'h0000005E: begin
				q			<=			16'h02C0;
		end
		32'h00000060: begin
				q			<=			16'hAA23;
		end
		32'h00000062: begin
				q			<=			16'h02D0;
		end
		32'h00000064: begin
				q			<=			16'hAC23;
		end
		32'h00000066: begin
				q			<=			16'h02E0;
		end
		32'h00000068: begin
				q			<=			16'hAE23;
		end
		32'h0000006A: begin
				q			<=			16'h02F0;
		end
		32'h0000006C: begin
				q			<=			16'hA023;
		end
		32'h0000006E: begin
				q			<=			16'h0500;
		end
		32'h00000070: begin
				q			<=			16'hA223;
		end
		32'h00000072: begin
				q			<=			16'h0510;
		end
		32'h00000074: begin
				q			<=			16'hA423;
		end
		32'h00000076: begin
				q			<=			16'h0520;
		end
		32'h00000078: begin
				q			<=			16'hA623;
		end
		32'h0000007A: begin
				q			<=			16'h0530;
		end
		32'h0000007C: begin
				q			<=			16'hA823;
		end
		32'h0000007E: begin
				q			<=			16'h0540;
		end
		32'h00000080: begin
				q			<=			16'hAA23;
		end
		32'h00000082: begin
				q			<=			16'h0550;
		end
		32'h00000084: begin
				q			<=			16'hAC23;
		end
		32'h00000086: begin
				q			<=			16'h0560;
		end
		32'h00000088: begin
				q			<=			16'hAE23;
		end
		32'h0000008A: begin
				q			<=			16'h0570;
		end
		32'h0000008C: begin
				q			<=			16'hA023;
		end
		32'h0000008E: begin
				q			<=			16'h0780;
		end
		32'h00000090: begin
				q			<=			16'hA223;
		end
		32'h00000092: begin
				q			<=			16'h0790;
		end
		32'h00000094: begin
				q			<=			16'hA423;
		end
		32'h00000096: begin
				q			<=			16'h07A0;
		end
		32'h00000098: begin
				q			<=			16'hA623;
		end
		32'h0000009A: begin
				q			<=			16'h07B0;
		end
		32'h0000009C: begin
				q			<=			16'hA823;
		end
		32'h0000009E: begin
				q			<=			16'h07C0;
		end
		32'h000000A0: begin
				q			<=			16'hAA23;
		end
		32'h000000A2: begin
				q			<=			16'h07D0;
		end
		32'h000000A4: begin
				q			<=			16'hAC23;
		end
		32'h000000A6: begin
				q			<=			16'h07E0;
		end
		32'h000000A8: begin
				q			<=			16'hAE23;
		end
		32'h000000AA: begin
				q			<=			16'h07F0;
		end
		32'h000000AC: begin
				q			<=			16'h0137;
		end
		32'h000000AE: begin
				q			<=			16'h0000;
		end
		32'h000000B0: begin
				q			<=			16'h0113;
		end
		32'h000000B2: begin
				q			<=			16'h3E01;
		end
		32'h000000B4: begin
				q			<=			16'h0537;
		end
		32'h000000B6: begin
				q			<=			16'h0000;
		end
		32'h000000B8: begin
				q			<=			16'h0513;
		end
		32'h000000BA: begin
				q			<=			16'h1605;
		end
		32'h000000BC: begin
				q			<=			16'hC58B;
		end
		32'h000000BE: begin
				q			<=			16'h0000;
		end
		32'h000000C0: begin
				q			<=			16'h00EF;
		end
		32'h000000C2: begin
				q			<=			16'h3FC0;
		end
		32'h000000C4: begin
				q			<=			16'h0093;
		end
		32'h000000C6: begin
				q			<=			16'h0005;
		end
		32'h000000C8: begin
				q			<=			16'hA103;
		end
		32'h000000CA: begin
				q			<=			16'h0000;
		end
		32'h000000CC: begin
				q			<=			16'h200B;
		end
		32'h000000CE: begin
				q			<=			16'h0201;
		end
		32'h000000D0: begin
				q			<=			16'hA103;
		end
		32'h000000D2: begin
				q			<=			16'h0040;
		end
		32'h000000D4: begin
				q			<=			16'h208B;
		end
		32'h000000D6: begin
				q			<=			16'h0201;
		end
		32'h000000D8: begin
				q			<=			16'hA103;
		end
		32'h000000DA: begin
				q			<=			16'h0080;
		end
		32'h000000DC: begin
				q			<=			16'h210B;
		end
		32'h000000DE: begin
				q			<=			16'h0201;
		end
		32'h000000E0: begin
				q			<=			16'hA183;
		end
		32'h000000E2: begin
				q			<=			16'h00C0;
		end
		32'h000000E4: begin
				q			<=			16'hA203;
		end
		32'h000000E6: begin
				q			<=			16'h0100;
		end
		32'h000000E8: begin
				q			<=			16'hA283;
		end
		32'h000000EA: begin
				q			<=			16'h0140;
		end
		32'h000000EC: begin
				q			<=			16'hA303;
		end
		32'h000000EE: begin
				q			<=			16'h0180;
		end
		32'h000000F0: begin
				q			<=			16'hA383;
		end
		32'h000000F2: begin
				q			<=			16'h01C0;
		end
		32'h000000F4: begin
				q			<=			16'hA403;
		end
		32'h000000F6: begin
				q			<=			16'h0200;
		end
		32'h000000F8: begin
				q			<=			16'hA483;
		end
		32'h000000FA: begin
				q			<=			16'h0240;
		end
		32'h000000FC: begin
				q			<=			16'hA503;
		end
		32'h000000FE: begin
				q			<=			16'h0280;
		end
		32'h00000100: begin
				q			<=			16'hA583;
		end
		32'h00000102: begin
				q			<=			16'h02C0;
		end
		32'h00000104: begin
				q			<=			16'hA603;
		end
		32'h00000106: begin
				q			<=			16'h0300;
		end
		32'h00000108: begin
				q			<=			16'hA683;
		end
		32'h0000010A: begin
				q			<=			16'h0340;
		end
		32'h0000010C: begin
				q			<=			16'hA703;
		end
		32'h0000010E: begin
				q			<=			16'h0380;
		end
		32'h00000110: begin
				q			<=			16'hA783;
		end
		32'h00000112: begin
				q			<=			16'h03C0;
		end
		32'h00000114: begin
				q			<=			16'hA803;
		end
		32'h00000116: begin
				q			<=			16'h0400;
		end
		32'h00000118: begin
				q			<=			16'hA883;
		end
		32'h0000011A: begin
				q			<=			16'h0440;
		end
		32'h0000011C: begin
				q			<=			16'hA903;
		end
		32'h0000011E: begin
				q			<=			16'h0480;
		end
		32'h00000120: begin
				q			<=			16'hA983;
		end
		32'h00000122: begin
				q			<=			16'h04C0;
		end
		32'h00000124: begin
				q			<=			16'hAA03;
		end
		32'h00000126: begin
				q			<=			16'h0500;
		end
		32'h00000128: begin
				q			<=			16'hAA83;
		end
		32'h0000012A: begin
				q			<=			16'h0540;
		end
		32'h0000012C: begin
				q			<=			16'hAB03;
		end
		32'h0000012E: begin
				q			<=			16'h0580;
		end
		32'h00000130: begin
				q			<=			16'hAB83;
		end
		32'h00000132: begin
				q			<=			16'h05C0;
		end
		32'h00000134: begin
				q			<=			16'hAC03;
		end
		32'h00000136: begin
				q			<=			16'h0600;
		end
		32'h00000138: begin
				q			<=			16'hAC83;
		end
		32'h0000013A: begin
				q			<=			16'h0640;
		end
		32'h0000013C: begin
				q			<=			16'hAD03;
		end
		32'h0000013E: begin
				q			<=			16'h0680;
		end
		32'h00000140: begin
				q			<=			16'hAD83;
		end
		32'h00000142: begin
				q			<=			16'h06C0;
		end
		32'h00000144: begin
				q			<=			16'hAE03;
		end
		32'h00000146: begin
				q			<=			16'h0700;
		end
		32'h00000148: begin
				q			<=			16'hAE83;
		end
		32'h0000014A: begin
				q			<=			16'h0740;
		end
		32'h0000014C: begin
				q			<=			16'hAF03;
		end
		32'h0000014E: begin
				q			<=			16'h0780;
		end
		32'h00000150: begin
				q			<=			16'hAF83;
		end
		32'h00000152: begin
				q			<=			16'h07C0;
		end
		32'h00000154: begin
				q			<=			16'hC08B;
		end
		32'h00000156: begin
				q			<=			16'h0000;
		end
		32'h00000158: begin
				q			<=			16'h410B;
		end
		32'h0000015A: begin
				q			<=			16'h0001;
		end
		32'h0000015C: begin
				q			<=			16'h000B;
		end
		32'h0000015E: begin
				q			<=			16'h0400;
		end
		32'h00000160: begin
				q			<=			16'h0000;
		end
		32'h00000162: begin
				q			<=			16'h0000;
		end
		32'h00000164: begin
				q			<=			16'h0000;
		end
		32'h00000166: begin
				q			<=			16'h0000;
		end
		32'h00000168: begin
				q			<=			16'h0000;
		end
		32'h0000016A: begin
				q			<=			16'h0000;
		end
		32'h0000016C: begin
				q			<=			16'h0000;
		end
		32'h0000016E: begin
				q			<=			16'h0000;
		end
		32'h00000170: begin
				q			<=			16'h0000;
		end
		32'h00000172: begin
				q			<=			16'h0000;
		end
		32'h00000174: begin
				q			<=			16'h0000;
		end
		32'h00000176: begin
				q			<=			16'h0000;
		end
		32'h00000178: begin
				q			<=			16'h0000;
		end
		32'h0000017A: begin
				q			<=			16'h0000;
		end
		32'h0000017C: begin
				q			<=			16'h0000;
		end
		32'h0000017E: begin
				q			<=			16'h0000;
		end
		32'h00000180: begin
				q			<=			16'h0000;
		end
		32'h00000182: begin
				q			<=			16'h0000;
		end
		32'h00000184: begin
				q			<=			16'h0000;
		end
		32'h00000186: begin
				q			<=			16'h0000;
		end
		32'h00000188: begin
				q			<=			16'h0000;
		end
		32'h0000018A: begin
				q			<=			16'h0000;
		end
		32'h0000018C: begin
				q			<=			16'h0000;
		end
		32'h0000018E: begin
				q			<=			16'h0000;
		end
		32'h00000190: begin
				q			<=			16'h0000;
		end
		32'h00000192: begin
				q			<=			16'h0000;
		end
		32'h00000194: begin
				q			<=			16'h0000;
		end
		32'h00000196: begin
				q			<=			16'h0000;
		end
		32'h00000198: begin
				q			<=			16'h0000;
		end
		32'h0000019A: begin
				q			<=			16'h0000;
		end
		32'h0000019C: begin
				q			<=			16'h0000;
		end
		32'h0000019E: begin
				q			<=			16'h0000;
		end
		32'h000001A0: begin
				q			<=			16'h0000;
		end
		32'h000001A2: begin
				q			<=			16'h0000;
		end
		32'h000001A4: begin
				q			<=			16'h0000;
		end
		32'h000001A6: begin
				q			<=			16'h0000;
		end
		32'h000001A8: begin
				q			<=			16'h0000;
		end
		32'h000001AA: begin
				q			<=			16'h0000;
		end
		32'h000001AC: begin
				q			<=			16'h0000;
		end
		32'h000001AE: begin
				q			<=			16'h0000;
		end
		32'h000001B0: begin
				q			<=			16'h0000;
		end
		32'h000001B2: begin
				q			<=			16'h0000;
		end
		32'h000001B4: begin
				q			<=			16'h0000;
		end
		32'h000001B6: begin
				q			<=			16'h0000;
		end
		32'h000001B8: begin
				q			<=			16'h0000;
		end
		32'h000001BA: begin
				q			<=			16'h0000;
		end
		32'h000001BC: begin
				q			<=			16'h0000;
		end
		32'h000001BE: begin
				q			<=			16'h0000;
		end
		32'h000001C0: begin
				q			<=			16'h0000;
		end
		32'h000001C2: begin
				q			<=			16'h0000;
		end
		32'h000001C4: begin
				q			<=			16'h0000;
		end
		32'h000001C6: begin
				q			<=			16'h0000;
		end
		32'h000001C8: begin
				q			<=			16'h0000;
		end
		32'h000001CA: begin
				q			<=			16'h0000;
		end
		32'h000001CC: begin
				q			<=			16'h0000;
		end
		32'h000001CE: begin
				q			<=			16'h0000;
		end
		32'h000001D0: begin
				q			<=			16'h0000;
		end
		32'h000001D2: begin
				q			<=			16'h0000;
		end
		32'h000001D4: begin
				q			<=			16'h0000;
		end
		32'h000001D6: begin
				q			<=			16'h0000;
		end
		32'h000001D8: begin
				q			<=			16'h0000;
		end
		32'h000001DA: begin
				q			<=			16'h0000;
		end
		32'h000001DC: begin
				q			<=			16'h0000;
		end
		32'h000001DE: begin
				q			<=			16'h0000;
		end
		32'h000001E0: begin
				q			<=			16'h0000;
		end
		32'h000001E2: begin
				q			<=			16'h0000;
		end
		32'h000001E4: begin
				q			<=			16'h0000;
		end
		32'h000001E6: begin
				q			<=			16'h0000;
		end
		32'h000001E8: begin
				q			<=			16'h0000;
		end
		32'h000001EA: begin
				q			<=			16'h0000;
		end
		32'h000001EC: begin
				q			<=			16'h0000;
		end
		32'h000001EE: begin
				q			<=			16'h0000;
		end
		32'h000001F0: begin
				q			<=			16'h0000;
		end
		32'h000001F2: begin
				q			<=			16'h0000;
		end
		32'h000001F4: begin
				q			<=			16'h0000;
		end
		32'h000001F6: begin
				q			<=			16'h0000;
		end
		32'h000001F8: begin
				q			<=			16'h0000;
		end
		32'h000001FA: begin
				q			<=			16'h0000;
		end
		32'h000001FC: begin
				q			<=			16'h0000;
		end
		32'h000001FE: begin
				q			<=			16'h0000;
		end
		32'h00000200: begin
				q			<=			16'h0000;
		end
		32'h00000202: begin
				q			<=			16'h0000;
		end
		32'h00000204: begin
				q			<=			16'h0000;
		end
		32'h00000206: begin
				q			<=			16'h0000;
		end
		32'h00000208: begin
				q			<=			16'h0000;
		end
		32'h0000020A: begin
				q			<=			16'h0000;
		end
		32'h0000020C: begin
				q			<=			16'h0000;
		end
		32'h0000020E: begin
				q			<=			16'h0000;
		end
		32'h00000210: begin
				q			<=			16'h0000;
		end
		32'h00000212: begin
				q			<=			16'h0000;
		end
		32'h00000214: begin
				q			<=			16'h0000;
		end
		32'h00000216: begin
				q			<=			16'h0000;
		end
		32'h00000218: begin
				q			<=			16'h0000;
		end
		32'h0000021A: begin
				q			<=			16'h0000;
		end
		32'h0000021C: begin
				q			<=			16'h0000;
		end
		32'h0000021E: begin
				q			<=			16'h0000;
		end
		32'h00000220: begin
				q			<=			16'h0000;
		end
		32'h00000222: begin
				q			<=			16'h0000;
		end
		32'h00000224: begin
				q			<=			16'h0000;
		end
		32'h00000226: begin
				q			<=			16'h0000;
		end
		32'h00000228: begin
				q			<=			16'h0000;
		end
		32'h0000022A: begin
				q			<=			16'h0000;
		end
		32'h0000022C: begin
				q			<=			16'h0000;
		end
		32'h0000022E: begin
				q			<=			16'h0000;
		end
		32'h00000230: begin
				q			<=			16'h0000;
		end
		32'h00000232: begin
				q			<=			16'h0000;
		end
		32'h00000234: begin
				q			<=			16'h0000;
		end
		32'h00000236: begin
				q			<=			16'h0000;
		end
		32'h00000238: begin
				q			<=			16'h0000;
		end
		32'h0000023A: begin
				q			<=			16'h0000;
		end
		32'h0000023C: begin
				q			<=			16'h0000;
		end
		32'h0000023E: begin
				q			<=			16'h0000;
		end
		32'h00000240: begin
				q			<=			16'h0000;
		end
		32'h00000242: begin
				q			<=			16'h0000;
		end
		32'h00000244: begin
				q			<=			16'h0000;
		end
		32'h00000246: begin
				q			<=			16'h0000;
		end
		32'h00000248: begin
				q			<=			16'h0000;
		end
		32'h0000024A: begin
				q			<=			16'h0000;
		end
		32'h0000024C: begin
				q			<=			16'h0000;
		end
		32'h0000024E: begin
				q			<=			16'h0000;
		end
		32'h00000250: begin
				q			<=			16'h0000;
		end
		32'h00000252: begin
				q			<=			16'h0000;
		end
		32'h00000254: begin
				q			<=			16'h0000;
		end
		32'h00000256: begin
				q			<=			16'h0000;
		end
		32'h00000258: begin
				q			<=			16'h0000;
		end
		32'h0000025A: begin
				q			<=			16'h0000;
		end
		32'h0000025C: begin
				q			<=			16'h0000;
		end
		32'h0000025E: begin
				q			<=			16'h0000;
		end
		32'h00000260: begin
				q			<=			16'h0000;
		end
		32'h00000262: begin
				q			<=			16'h0000;
		end
		32'h00000264: begin
				q			<=			16'h0000;
		end
		32'h00000266: begin
				q			<=			16'h0000;
		end
		32'h00000268: begin
				q			<=			16'h0000;
		end
		32'h0000026A: begin
				q			<=			16'h0000;
		end
		32'h0000026C: begin
				q			<=			16'h0000;
		end
		32'h0000026E: begin
				q			<=			16'h0000;
		end
		32'h00000270: begin
				q			<=			16'h0000;
		end
		32'h00000272: begin
				q			<=			16'h0000;
		end
		32'h00000274: begin
				q			<=			16'h0000;
		end
		32'h00000276: begin
				q			<=			16'h0000;
		end
		32'h00000278: begin
				q			<=			16'h0000;
		end
		32'h0000027A: begin
				q			<=			16'h0000;
		end
		32'h0000027C: begin
				q			<=			16'h0000;
		end
		32'h0000027E: begin
				q			<=			16'h0000;
		end
		32'h00000280: begin
				q			<=			16'h0000;
		end
		32'h00000282: begin
				q			<=			16'h0000;
		end
		32'h00000284: begin
				q			<=			16'h0000;
		end
		32'h00000286: begin
				q			<=			16'h0000;
		end
		32'h00000288: begin
				q			<=			16'h0000;
		end
		32'h0000028A: begin
				q			<=			16'h0000;
		end
		32'h0000028C: begin
				q			<=			16'h0000;
		end
		32'h0000028E: begin
				q			<=			16'h0000;
		end
		32'h00000290: begin
				q			<=			16'h0000;
		end
		32'h00000292: begin
				q			<=			16'h0000;
		end
		32'h00000294: begin
				q			<=			16'h0000;
		end
		32'h00000296: begin
				q			<=			16'h0000;
		end
		32'h00000298: begin
				q			<=			16'h0000;
		end
		32'h0000029A: begin
				q			<=			16'h0000;
		end
		32'h0000029C: begin
				q			<=			16'h0000;
		end
		32'h0000029E: begin
				q			<=			16'h0000;
		end
		32'h000002A0: begin
				q			<=			16'h0000;
		end
		32'h000002A2: begin
				q			<=			16'h0000;
		end
		32'h000002A4: begin
				q			<=			16'h0000;
		end
		32'h000002A6: begin
				q			<=			16'h0000;
		end
		32'h000002A8: begin
				q			<=			16'h0000;
		end
		32'h000002AA: begin
				q			<=			16'h0000;
		end
		32'h000002AC: begin
				q			<=			16'h0000;
		end
		32'h000002AE: begin
				q			<=			16'h0000;
		end
		32'h000002B0: begin
				q			<=			16'h0000;
		end
		32'h000002B2: begin
				q			<=			16'h0000;
		end
		32'h000002B4: begin
				q			<=			16'h0000;
		end
		32'h000002B6: begin
				q			<=			16'h0000;
		end
		32'h000002B8: begin
				q			<=			16'h0000;
		end
		32'h000002BA: begin
				q			<=			16'h0000;
		end
		32'h000002BC: begin
				q			<=			16'h0000;
		end
		32'h000002BE: begin
				q			<=			16'h0000;
		end
		32'h000002C0: begin
				q			<=			16'h0000;
		end
		32'h000002C2: begin
				q			<=			16'h0000;
		end
		32'h000002C4: begin
				q			<=			16'h0000;
		end
		32'h000002C6: begin
				q			<=			16'h0000;
		end
		32'h000002C8: begin
				q			<=			16'h0000;
		end
		32'h000002CA: begin
				q			<=			16'h0000;
		end
		32'h000002CC: begin
				q			<=			16'h0000;
		end
		32'h000002CE: begin
				q			<=			16'h0000;
		end
		32'h000002D0: begin
				q			<=			16'h0000;
		end
		32'h000002D2: begin
				q			<=			16'h0000;
		end
		32'h000002D4: begin
				q			<=			16'h0000;
		end
		32'h000002D6: begin
				q			<=			16'h0000;
		end
		32'h000002D8: begin
				q			<=			16'h0000;
		end
		32'h000002DA: begin
				q			<=			16'h0000;
		end
		32'h000002DC: begin
				q			<=			16'h0000;
		end
		32'h000002DE: begin
				q			<=			16'h0000;
		end
		32'h000002E0: begin
				q			<=			16'h0000;
		end
		32'h000002E2: begin
				q			<=			16'h0000;
		end
		32'h000002E4: begin
				q			<=			16'h0000;
		end
		32'h000002E6: begin
				q			<=			16'h0000;
		end
		32'h000002E8: begin
				q			<=			16'h0000;
		end
		32'h000002EA: begin
				q			<=			16'h0000;
		end
		32'h000002EC: begin
				q			<=			16'h0000;
		end
		32'h000002EE: begin
				q			<=			16'h0000;
		end
		32'h000002F0: begin
				q			<=			16'h0000;
		end
		32'h000002F2: begin
				q			<=			16'h0000;
		end
		32'h000002F4: begin
				q			<=			16'h0000;
		end
		32'h000002F6: begin
				q			<=			16'h0000;
		end
		32'h000002F8: begin
				q			<=			16'h0000;
		end
		32'h000002FA: begin
				q			<=			16'h0000;
		end
		32'h000002FC: begin
				q			<=			16'h0000;
		end
		32'h000002FE: begin
				q			<=			16'h0000;
		end
		32'h00000300: begin
				q			<=			16'h0000;
		end
		32'h00000302: begin
				q			<=			16'h0000;
		end
		32'h00000304: begin
				q			<=			16'h0000;
		end
		32'h00000306: begin
				q			<=			16'h0000;
		end
		32'h00000308: begin
				q			<=			16'h0000;
		end
		32'h0000030A: begin
				q			<=			16'h0000;
		end
		32'h0000030C: begin
				q			<=			16'h0000;
		end
		32'h0000030E: begin
				q			<=			16'h0000;
		end
		32'h00000310: begin
				q			<=			16'h0000;
		end
		32'h00000312: begin
				q			<=			16'h0000;
		end
		32'h00000314: begin
				q			<=			16'h0000;
		end
		32'h00000316: begin
				q			<=			16'h0000;
		end
		32'h00000318: begin
				q			<=			16'h0000;
		end
		32'h0000031A: begin
				q			<=			16'h0000;
		end
		32'h0000031C: begin
				q			<=			16'h0000;
		end
		32'h0000031E: begin
				q			<=			16'h0000;
		end
		32'h00000320: begin
				q			<=			16'h0000;
		end
		32'h00000322: begin
				q			<=			16'h0000;
		end
		32'h00000324: begin
				q			<=			16'h0000;
		end
		32'h00000326: begin
				q			<=			16'h0000;
		end
		32'h00000328: begin
				q			<=			16'h0000;
		end
		32'h0000032A: begin
				q			<=			16'h0000;
		end
		32'h0000032C: begin
				q			<=			16'h0000;
		end
		32'h0000032E: begin
				q			<=			16'h0000;
		end
		32'h00000330: begin
				q			<=			16'h0000;
		end
		32'h00000332: begin
				q			<=			16'h0000;
		end
		32'h00000334: begin
				q			<=			16'h0000;
		end
		32'h00000336: begin
				q			<=			16'h0000;
		end
		32'h00000338: begin
				q			<=			16'h0000;
		end
		32'h0000033A: begin
				q			<=			16'h0000;
		end
		32'h0000033C: begin
				q			<=			16'h0000;
		end
		32'h0000033E: begin
				q			<=			16'h0000;
		end
		32'h00000340: begin
				q			<=			16'h0000;
		end
		32'h00000342: begin
				q			<=			16'h0000;
		end
		32'h00000344: begin
				q			<=			16'h0000;
		end
		32'h00000346: begin
				q			<=			16'h0000;
		end
		32'h00000348: begin
				q			<=			16'h0000;
		end
		32'h0000034A: begin
				q			<=			16'h0000;
		end
		32'h0000034C: begin
				q			<=			16'h0000;
		end
		32'h0000034E: begin
				q			<=			16'h0000;
		end
		32'h00000350: begin
				q			<=			16'h0000;
		end
		32'h00000352: begin
				q			<=			16'h0000;
		end
		32'h00000354: begin
				q			<=			16'h0000;
		end
		32'h00000356: begin
				q			<=			16'h0000;
		end
		32'h00000358: begin
				q			<=			16'h0000;
		end
		32'h0000035A: begin
				q			<=			16'h0000;
		end
		32'h0000035C: begin
				q			<=			16'h0000;
		end
		32'h0000035E: begin
				q			<=			16'h0000;
		end
		32'h00000360: begin
				q			<=			16'h0000;
		end
		32'h00000362: begin
				q			<=			16'h0000;
		end
		32'h00000364: begin
				q			<=			16'h0000;
		end
		32'h00000366: begin
				q			<=			16'h0000;
		end
		32'h00000368: begin
				q			<=			16'h0000;
		end
		32'h0000036A: begin
				q			<=			16'h0000;
		end
		32'h0000036C: begin
				q			<=			16'h0000;
		end
		32'h0000036E: begin
				q			<=			16'h0000;
		end
		32'h00000370: begin
				q			<=			16'h0000;
		end
		32'h00000372: begin
				q			<=			16'h0000;
		end
		32'h00000374: begin
				q			<=			16'h0000;
		end
		32'h00000376: begin
				q			<=			16'h0000;
		end
		32'h00000378: begin
				q			<=			16'h0000;
		end
		32'h0000037A: begin
				q			<=			16'h0000;
		end
		32'h0000037C: begin
				q			<=			16'h0000;
		end
		32'h0000037E: begin
				q			<=			16'h0000;
		end
		32'h00000380: begin
				q			<=			16'h0000;
		end
		32'h00000382: begin
				q			<=			16'h0000;
		end
		32'h00000384: begin
				q			<=			16'h0000;
		end
		32'h00000386: begin
				q			<=			16'h0000;
		end
		32'h00000388: begin
				q			<=			16'h0000;
		end
		32'h0000038A: begin
				q			<=			16'h0000;
		end
		32'h0000038C: begin
				q			<=			16'h0000;
		end
		32'h0000038E: begin
				q			<=			16'h0000;
		end
		32'h00000390: begin
				q			<=			16'h0000;
		end
		32'h00000392: begin
				q			<=			16'h0000;
		end
		32'h00000394: begin
				q			<=			16'h0000;
		end
		32'h00000396: begin
				q			<=			16'h0000;
		end
		32'h00000398: begin
				q			<=			16'h0000;
		end
		32'h0000039A: begin
				q			<=			16'h0000;
		end
		32'h0000039C: begin
				q			<=			16'h0000;
		end
		32'h0000039E: begin
				q			<=			16'h0000;
		end
		32'h000003A0: begin
				q			<=			16'h0000;
		end
		32'h000003A2: begin
				q			<=			16'h0000;
		end
		32'h000003A4: begin
				q			<=			16'h0000;
		end
		32'h000003A6: begin
				q			<=			16'h0000;
		end
		32'h000003A8: begin
				q			<=			16'h0000;
		end
		32'h000003AA: begin
				q			<=			16'h0000;
		end
		32'h000003AC: begin
				q			<=			16'h0000;
		end
		32'h000003AE: begin
				q			<=			16'h0000;
		end
		32'h000003B0: begin
				q			<=			16'h0000;
		end
		32'h000003B2: begin
				q			<=			16'h0000;
		end
		32'h000003B4: begin
				q			<=			16'h0000;
		end
		32'h000003B6: begin
				q			<=			16'h0000;
		end
		32'h000003B8: begin
				q			<=			16'h0000;
		end
		32'h000003BA: begin
				q			<=			16'h0000;
		end
		32'h000003BC: begin
				q			<=			16'h0000;
		end
		32'h000003BE: begin
				q			<=			16'h0000;
		end
		32'h000003C0: begin
				q			<=			16'h0000;
		end
		32'h000003C2: begin
				q			<=			16'h0000;
		end
		32'h000003C4: begin
				q			<=			16'h0000;
		end
		32'h000003C6: begin
				q			<=			16'h0000;
		end
		32'h000003C8: begin
				q			<=			16'h0000;
		end
		32'h000003CA: begin
				q			<=			16'h0000;
		end
		32'h000003CC: begin
				q			<=			16'h0000;
		end
		32'h000003CE: begin
				q			<=			16'h0000;
		end
		32'h000003D0: begin
				q			<=			16'h0000;
		end
		32'h000003D2: begin
				q			<=			16'h0000;
		end
		32'h000003D4: begin
				q			<=			16'h0000;
		end
		32'h000003D6: begin
				q			<=			16'h0000;
		end
		32'h000003D8: begin
				q			<=			16'h0000;
		end
		32'h000003DA: begin
				q			<=			16'h0000;
		end
		32'h000003DC: begin
				q			<=			16'h0000;
		end
		32'h000003DE: begin
				q			<=			16'h0000;
		end
		32'h000003E0: begin
				q			<=			16'h00EF;
		end
		32'h000003E2: begin
				q			<=			16'h0180;
		end
		32'h000003E4: begin
				q			<=			16'h0073;
		end
		32'h000003E6: begin
				q			<=			16'h0010;
		end
		32'h000003E8: begin
				q			<=			16'h0000;
		end
		32'h000003EA: begin
				q			<=			16'h0000;
		end
		32'h000003EC: begin
				q			<=			16'h0000;
		end
		32'h000003EE: begin
				q			<=			16'h0000;
		end
		32'h000003F0: begin
				q			<=			16'h0000;
		end
		32'h000003F2: begin
				q			<=			16'h0000;
		end
		32'h000003F4: begin
				q			<=			16'h0000;
		end
		32'h000003F6: begin
				q			<=			16'h0000;
		end
		32'h000003F8: begin
				q			<=			16'h0113;
		end
		32'h000003FA: begin
				q			<=			16'hFF01;
		end
		32'h000003FC: begin
				q			<=			16'h2623;
		end
		32'h000003FE: begin
				q			<=			16'h0011;
		end
		32'h00000400: begin
				q			<=			16'h17B7;
		end
		32'h00000402: begin
				q			<=			16'h0001;
		end
		32'h00000404: begin
				q			<=			16'h8C23;
		end
		32'h00000406: begin
				q			<=			16'hF807;
		end
		32'h00000408: begin
				q			<=			16'h1737;
		end
		32'h0000040A: begin
				q			<=			16'h0001;
		end
		32'h0000040C: begin
				q			<=			16'h0713;
		end
		32'h0000040E: begin
				q			<=			16'h8F47;
		end
		32'h00000410: begin
				q			<=			16'h17B7;
		end
		32'h00000412: begin
				q			<=			16'h0001;
		end
		32'h00000414: begin
				q			<=			16'h8793;
		end
		32'h00000416: begin
				q			<=			16'hF707;
		end
		32'h00000418: begin
				q			<=			16'h7063;
		end
		32'h0000041A: begin
				q			<=			16'h02F7;
		end
		32'h0000041C: begin
				q			<=			16'h17B7;
		end
		32'h0000041E: begin
				q			<=			16'h0001;
		end
		32'h00000420: begin
				q			<=			16'h8793;
		end
		32'h00000422: begin
				q			<=			16'h8F47;
		end
		32'h00000424: begin
				q			<=			16'h1737;
		end
		32'h00000426: begin
				q			<=			16'h0001;
		end
		32'h00000428: begin
				q			<=			16'h0713;
		end
		32'h0000042A: begin
				q			<=			16'hF707;
		end
		32'h0000042C: begin
				q			<=			16'hA023;
		end
		32'h0000042E: begin
				q			<=			16'h0007;
		end
		32'h00000430: begin
				q			<=			16'h8793;
		end
		32'h00000432: begin
				q			<=			16'h0047;
		end
		32'h00000434: begin
				q			<=			16'hECE3;
		end
		32'h00000436: begin
				q			<=			16'hFEE7;
		end
		32'h00000438: begin
				q			<=			16'h0513;
		end
		32'h0000043A: begin
				q			<=			16'h0000;
		end
		32'h0000043C: begin
				q			<=			16'h00EF;
		end
		32'h0000043E: begin
				q			<=			16'h6550;
		end
		32'h00000440: begin
				q			<=			16'h00EF;
		end
		32'h00000442: begin
				q			<=			16'h0140;
		end
		32'h00000444: begin
				q			<=			16'h2083;
		end
		32'h00000446: begin
				q			<=			16'h00C1;
		end
		32'h00000448: begin
				q			<=			16'h0113;
		end
		32'h0000044A: begin
				q			<=			16'h0101;
		end
		32'h0000044C: begin
				q			<=			16'h8067;
		end
		32'h0000044E: begin
				q			<=			16'h0000;
		end
		32'h00000450: begin
				q			<=			16'h0000;
		end
		32'h00000452: begin
				q			<=			16'h0000;
		end
		32'h00000454: begin
				q			<=			16'h0113;
		end
		32'h00000456: begin
				q			<=			16'hFF01;
		end
		32'h00000458: begin
				q			<=			16'h2623;
		end
		32'h0000045A: begin
				q			<=			16'h0011;
		end
		32'h0000045C: begin
				q			<=			16'h2423;
		end
		32'h0000045E: begin
				q			<=			16'h0081;
		end
		32'h00000460: begin
				q			<=			16'h0513;
		end
		32'h00000462: begin
				q			<=			16'h0000;
		end
		32'h00000464: begin
				q			<=			16'h00EF;
		end
		32'h00000466: begin
				q			<=			16'h0EC0;
		end
		32'h00000468: begin
				q			<=			16'h0537;
		end
		32'h0000046A: begin
				q			<=			16'h0100;
		end
		32'h0000046C: begin
				q			<=			16'h00EF;
		end
		32'h0000046E: begin
				q			<=			16'h0F80;
		end
		32'h00000470: begin
				q			<=			16'h0537;
		end
		32'h00000472: begin
				q			<=			16'h0180;
		end
		32'h00000474: begin
				q			<=			16'h00EF;
		end
		32'h00000476: begin
				q			<=			16'h1080;
		end
		32'h00000478: begin
				q			<=			16'h00EF;
		end
		32'h0000047A: begin
				q			<=			16'h11C0;
		end
		32'h0000047C: begin
				q			<=			16'h17B7;
		end
		32'h0000047E: begin
				q			<=			16'h0001;
		end
		32'h00000480: begin
				q			<=			16'h0713;
		end
		32'h00000482: begin
				q			<=			16'h0010;
		end
		32'h00000484: begin
				q			<=			16'h8C23;
		end
		32'h00000486: begin
				q			<=			16'hF8E7;
		end
		32'h00000488: begin
				q			<=			16'h00EF;
		end
		32'h0000048A: begin
				q			<=			16'h1480;
		end
		32'h0000048C: begin
				q			<=			16'h5437;
		end
		32'h0000048E: begin
				q			<=			16'h0000;
		end
		32'h00000490: begin
				q			<=			16'h006F;
		end
		32'h00000492: begin
				q			<=			16'h0080;
		end
		32'h00000494: begin
				q			<=			16'h00EF;
		end
		32'h00000496: begin
				q			<=			16'h1280;
		end
		32'h00000498: begin
				q			<=			16'h0793;
		end
		32'h0000049A: begin
				q			<=			16'hE204;
		end
		32'h0000049C: begin
				q			<=			16'h8793;
		end
		32'h0000049E: begin
				q			<=			16'hFFF7;
		end
		32'h000004A0: begin
				q			<=			16'h9EE3;
		end
		32'h000004A2: begin
				q			<=			16'hFE07;
		end
		32'h000004A4: begin
				q			<=			16'hF06F;
		end
		32'h000004A6: begin
				q			<=			16'hFF1F;
		end
		32'h000004A8: begin
				q			<=			16'h0000;
		end
		32'h000004AA: begin
				q			<=			16'h0000;
		end
		32'h000004AC: begin
				q			<=			16'h07B7;
		end
		32'h000004AE: begin
				q			<=			16'h8000;
		end
		32'h000004B0: begin
				q			<=			16'hA503;
		end
		32'h000004B2: begin
				q			<=			16'h0107;
		end
		32'h000004B4: begin
				q			<=			16'h8067;
		end
		32'h000004B6: begin
				q			<=			16'h0000;
		end
		32'h000004B8: begin
				q			<=			16'h0000;
		end
		32'h000004BA: begin
				q			<=			16'h0000;
		end
		32'h000004BC: begin
				q			<=			16'h0113;
		end
		32'h000004BE: begin
				q			<=			16'hFF01;
		end
		32'h000004C0: begin
				q			<=			16'h2623;
		end
		32'h000004C2: begin
				q			<=			16'h0011;
		end
		32'h000004C4: begin
				q			<=			16'h2423;
		end
		32'h000004C6: begin
				q			<=			16'h0081;
		end
		32'h000004C8: begin
				q			<=			16'h2223;
		end
		32'h000004CA: begin
				q			<=			16'h0091;
		end
		32'h000004CC: begin
				q			<=			16'h0493;
		end
		32'h000004CE: begin
				q			<=			16'h0005;
		end
		32'h000004D0: begin
				q			<=			16'h17B7;
		end
		32'h000004D2: begin
				q			<=			16'h0001;
		end
		32'h000004D4: begin
				q			<=			16'hC783;
		end
		32'h000004D6: begin
				q			<=			16'hF987;
		end
		32'h000004D8: begin
				q			<=			16'h8463;
		end
		32'h000004DA: begin
				q			<=			16'h0207;
		end
		32'h000004DC: begin
				q			<=			16'h8413;
		end
		32'h000004DE: begin
				q			<=			16'h0005;
		end
		32'h000004E0: begin
				q			<=			16'hF793;
		end
		32'h000004E2: begin
				q			<=			16'h0085;
		end
		32'h000004E4: begin
				q			<=			16'h8A63;
		end
		32'h000004E6: begin
				q			<=			16'h0007;
		end
		32'h000004E8: begin
				q			<=			16'h17B7;
		end
		32'h000004EA: begin
				q			<=			16'h0001;
		end
		32'h000004EC: begin
				q			<=			16'hA703;
		end
		32'h000004EE: begin
				q			<=			16'hF747;
		end
		32'h000004F0: begin
				q			<=			16'h0793;
		end
		32'h000004F2: begin
				q			<=			16'h0010;
		end
		32'h000004F4: begin
				q			<=			16'h0263;
		end
		32'h000004F6: begin
				q			<=			16'h02F7;
		end
		32'h000004F8: begin
				q			<=			16'h7413;
		end
		32'h000004FA: begin
				q			<=			16'h0104;
		end
		32'h000004FC: begin
				q			<=			16'h1E63;
		end
		32'h000004FE: begin
				q			<=			16'h0204;
		end
		32'h00000500: begin
				q			<=			16'h8513;
		end
		32'h00000502: begin
				q			<=			16'h0004;
		end
		32'h00000504: begin
				q			<=			16'h2083;
		end
		32'h00000506: begin
				q			<=			16'h00C1;
		end
		32'h00000508: begin
				q			<=			16'h2403;
		end
		32'h0000050A: begin
				q			<=			16'h0081;
		end
		32'h0000050C: begin
				q			<=			16'h2483;
		end
		32'h0000050E: begin
				q			<=			16'h0041;
		end
		32'h00000510: begin
				q			<=			16'h0113;
		end
		32'h00000512: begin
				q			<=			16'h0101;
		end
		32'h00000514: begin
				q			<=			16'h8067;
		end
		32'h00000516: begin
				q			<=			16'h0000;
		end
		32'h00000518: begin
				q			<=			16'h17B7;
		end
		32'h0000051A: begin
				q			<=			16'h0001;
		end
		32'h0000051C: begin
				q			<=			16'hA703;
		end
		32'h0000051E: begin
				q			<=			16'hF847;
		end
		32'h00000520: begin
				q			<=			16'h0793;
		end
		32'h00000522: begin
				q			<=			16'h0010;
		end
		32'h00000524: begin
				q			<=			16'h1AE3;
		end
		32'h00000526: begin
				q			<=			16'hFCF7;
		end
		32'h00000528: begin
				q			<=			16'h17B7;
		end
		32'h0000052A: begin
				q			<=			16'h0001;
		end
		32'h0000052C: begin
				q			<=			16'hA223;
		end
		32'h0000052E: begin
				q			<=			16'hF807;
		end
		32'h00000530: begin
				q			<=			16'h00EF;
		end
		32'h00000532: begin
				q			<=			16'h0640;
		end
		32'h00000534: begin
				q			<=			16'hF06F;
		end
		32'h00000536: begin
				q			<=			16'hFC5F;
		end
		32'h00000538: begin
				q			<=			16'h07B7;
		end
		32'h0000053A: begin
				q			<=			16'h8000;
		end
		32'h0000053C: begin
				q			<=			16'hA503;
		end
		32'h0000053E: begin
				q			<=			16'h0207;
		end
		32'h00000540: begin
				q			<=			16'h7513;
		end
		32'h00000542: begin
				q			<=			16'h0FF5;
		end
		32'h00000544: begin
				q			<=			16'h00EF;
		end
		32'h00000546: begin
				q			<=			16'h5940;
		end
		32'h00000548: begin
				q			<=			16'hF06F;
		end
		32'h0000054A: begin
				q			<=			16'hFB9F;
		end
		32'h0000054C: begin
				q			<=			16'h0000;
		end
		32'h0000054E: begin
				q			<=			16'h0000;
		end
		32'h00000550: begin
				q			<=			16'h7513;
		end
		32'h00000552: begin
				q			<=			16'h01F5;
		end
		32'h00000554: begin
				q			<=			16'h07B7;
		end
		32'h00000556: begin
				q			<=			16'h8000;
		end
		32'h00000558: begin
				q			<=			16'hA423;
		end
		32'h0000055A: begin
				q			<=			16'h02A7;
		end
		32'h0000055C: begin
				q			<=			16'h8067;
		end
		32'h0000055E: begin
				q			<=			16'h0000;
		end
		32'h00000560: begin
				q			<=			16'h0000;
		end
		32'h00000562: begin
				q			<=			16'h0000;
		end
		32'h00000564: begin
				q			<=			16'h17B7;
		end
		32'h00000566: begin
				q			<=			16'h0001;
		end
		32'h00000568: begin
				q			<=			16'hAE23;
		end
		32'h0000056A: begin
				q			<=			16'hF6A7;
		end
		32'h0000056C: begin
				q			<=			16'h07B7;
		end
		32'h0000056E: begin
				q			<=			16'h8000;
		end
		32'h00000570: begin
				q			<=			16'hA823;
		end
		32'h00000572: begin
				q			<=			16'h02A7;
		end
		32'h00000574: begin
				q			<=			16'h8067;
		end
		32'h00000576: begin
				q			<=			16'h0000;
		end
		32'h00000578: begin
				q			<=			16'h0000;
		end
		32'h0000057A: begin
				q			<=			16'h0000;
		end
		32'h0000057C: begin
				q			<=			16'h17B7;
		end
		32'h0000057E: begin
				q			<=			16'h0001;
		end
		32'h00000580: begin
				q			<=			16'hA023;
		end
		32'h00000582: begin
				q			<=			16'hF8A7;
		end
		32'h00000584: begin
				q			<=			16'h07B7;
		end
		32'h00000586: begin
				q			<=			16'h8000;
		end
		32'h00000588: begin
				q			<=			16'hAA23;
		end
		32'h0000058A: begin
				q			<=			16'h02A7;
		end
		32'h0000058C: begin
				q			<=			16'h8067;
		end
		32'h0000058E: begin
				q			<=			16'h0000;
		end
		32'h00000590: begin
				q			<=			16'h0000;
		end
		32'h00000592: begin
				q			<=			16'h0000;
		end
		32'h00000594: begin
				q			<=			16'h07B7;
		end
		32'h00000596: begin
				q			<=			16'h8000;
		end
		32'h00000598: begin
				q			<=			16'h0713;
		end
		32'h0000059A: begin
				q			<=			16'h0010;
		end
		32'h0000059C: begin
				q			<=			16'hA623;
		end
		32'h0000059E: begin
				q			<=			16'h02E7;
		end
		32'h000005A0: begin
				q			<=			16'h17B7;
		end
		32'h000005A2: begin
				q			<=			16'h0001;
		end
		32'h000005A4: begin
				q			<=			16'h8793;
		end
		32'h000005A6: begin
				q			<=			16'hF787;
		end
		32'h000005A8: begin
				q			<=			16'hA703;
		end
		32'h000005AA: begin
				q			<=			16'h0007;
		end
		32'h000005AC: begin
				q			<=			16'h3713;
		end
		32'h000005AE: begin
				q			<=			16'h0017;
		end
		32'h000005B0: begin
				q			<=			16'hA023;
		end
		32'h000005B2: begin
				q			<=			16'h00E7;
		end
		32'h000005B4: begin
				q			<=			16'h8067;
		end
		32'h000005B6: begin
				q			<=			16'h0000;
		end
		32'h000005B8: begin
				q			<=			16'h0000;
		end
		32'h000005BA: begin
				q			<=			16'h0000;
		end
		32'h000005BC: begin
				q			<=			16'h17B7;
		end
		32'h000005BE: begin
				q			<=			16'h0001;
		end
		32'h000005C0: begin
				q			<=			16'h0713;
		end
		32'h000005C2: begin
				q			<=			16'h0010;
		end
		32'h000005C4: begin
				q			<=			16'hA223;
		end
		32'h000005C6: begin
				q			<=			16'hF8E7;
		end
		32'h000005C8: begin
				q			<=			16'h8067;
		end
		32'h000005CA: begin
				q			<=			16'h0000;
		end
		32'h000005CC: begin
				q			<=			16'h0000;
		end
		32'h000005CE: begin
				q			<=			16'h0000;
		end
		32'h000005D0: begin
				q			<=			16'h17B7;
		end
		32'h000005D2: begin
				q			<=			16'h0001;
		end
		32'h000005D4: begin
				q			<=			16'h0713;
		end
		32'h000005D6: begin
				q			<=			16'h0010;
		end
		32'h000005D8: begin
				q			<=			16'hAA23;
		end
		32'h000005DA: begin
				q			<=			16'hF6E7;
		end
		32'h000005DC: begin
				q			<=			16'h8067;
		end
		32'h000005DE: begin
				q			<=			16'h0000;
		end
		32'h000005E0: begin
				q			<=			16'h0000;
		end
		32'h000005E2: begin
				q			<=			16'h0000;
		end
		32'h000005E4: begin
				q			<=			16'h17B7;
		end
		32'h000005E6: begin
				q			<=			16'h0001;
		end
		32'h000005E8: begin
				q			<=			16'hAA23;
		end
		32'h000005EA: begin
				q			<=			16'hF607;
		end
		32'h000005EC: begin
				q			<=			16'h8067;
		end
		32'h000005EE: begin
				q			<=			16'h0000;
		end
		32'h000005F0: begin
				q			<=			16'h0000;
		end
		32'h000005F2: begin
				q			<=			16'h0000;
		end
		32'h000005F4: begin
				q			<=			16'h17B7;
		end
		32'h000005F6: begin
				q			<=			16'h0001;
		end
		32'h000005F8: begin
				q			<=			16'hA783;
		end
		32'h000005FA: begin
				q			<=			16'hF787;
		end
		32'h000005FC: begin
				q			<=			16'h8863;
		end
		32'h000005FE: begin
				q			<=			16'h0007;
		end
		32'h00000600: begin
				q			<=			16'h0713;
		end
		32'h00000602: begin
				q			<=			16'h0010;
		end
		32'h00000604: begin
				q			<=			16'h8263;
		end
		32'h00000606: begin
				q			<=			16'h02E7;
		end
		32'h00000608: begin
				q			<=			16'h8067;
		end
		32'h0000060A: begin
				q			<=			16'h0000;
		end
		32'h0000060C: begin
				q			<=			16'h17B7;
		end
		32'h0000060E: begin
				q			<=			16'h0001;
		end
		32'h00000610: begin
				q			<=			16'hA783;
		end
		32'h00000612: begin
				q			<=			16'hF807;
		end
		32'h00000614: begin
				q			<=			16'h0533;
		end
		32'h00000616: begin
				q			<=			16'h00F5;
		end
		32'h00000618: begin
				q			<=			16'h07B7;
		end
		32'h0000061A: begin
				q			<=			16'h4000;
		end
		32'h0000061C: begin
				q			<=			16'h6533;
		end
		32'h0000061E: begin
				q			<=			16'h00F5;
		end
		32'h00000620: begin
				q			<=			16'h2023;
		end
		32'h00000622: begin
				q			<=			16'h00B5;
		end
		32'h00000624: begin
				q			<=			16'h8067;
		end
		32'h00000626: begin
				q			<=			16'h0000;
		end
		32'h00000628: begin
				q			<=			16'h17B7;
		end
		32'h0000062A: begin
				q			<=			16'h0001;
		end
		32'h0000062C: begin
				q			<=			16'hA783;
		end
		32'h0000062E: begin
				q			<=			16'hF7C7;
		end
		32'h00000630: begin
				q			<=			16'h0533;
		end
		32'h00000632: begin
				q			<=			16'h00F5;
		end
		32'h00000634: begin
				q			<=			16'h07B7;
		end
		32'h00000636: begin
				q			<=			16'h4000;
		end
		32'h00000638: begin
				q			<=			16'h6533;
		end
		32'h0000063A: begin
				q			<=			16'h00F5;
		end
		32'h0000063C: begin
				q			<=			16'h2023;
		end
		32'h0000063E: begin
				q			<=			16'h00B5;
		end
		32'h00000640: begin
				q			<=			16'hF06F;
		end
		32'h00000642: begin
				q			<=			16'hFC9F;
		end
		32'h00000644: begin
				q			<=			16'h0000;
		end
		32'h00000646: begin
				q			<=			16'h0000;
		end
		32'h00000648: begin
				q			<=			16'h17B7;
		end
		32'h0000064A: begin
				q			<=			16'h0001;
		end
		32'h0000064C: begin
				q			<=			16'hA783;
		end
		32'h0000064E: begin
				q			<=			16'hF787;
		end
		32'h00000650: begin
				q			<=			16'h9863;
		end
		32'h00000652: begin
				q			<=			16'h0207;
		end
		32'h00000654: begin
				q			<=			16'h0713;
		end
		32'h00000656: begin
				q			<=			16'h0000;
		end
		32'h00000658: begin
				q			<=			16'h15B7;
		end
		32'h0000065A: begin
				q			<=			16'h0001;
		end
		32'h0000065C: begin
				q			<=			16'h0637;
		end
		32'h0000065E: begin
				q			<=			16'h4000;
		end
		32'h00000660: begin
				q			<=			16'h66B7;
		end
		32'h00000662: begin
				q			<=			16'h0009;
		end
		32'h00000664: begin
				q			<=			16'hA783;
		end
		32'h00000666: begin
				q			<=			16'hF805;
		end
		32'h00000668: begin
				q			<=			16'h07B3;
		end
		32'h0000066A: begin
				q			<=			16'h00F7;
		end
		32'h0000066C: begin
				q			<=			16'hE7B3;
		end
		32'h0000066E: begin
				q			<=			16'h00C7;
		end
		32'h00000670: begin
				q			<=			16'hA023;
		end
		32'h00000672: begin
				q			<=			16'h0007;
		end
		32'h00000674: begin
				q			<=			16'h0713;
		end
		32'h00000676: begin
				q			<=			16'h0047;
		end
		32'h00000678: begin
				q			<=			16'h16E3;
		end
		32'h0000067A: begin
				q			<=			16'hFED7;
		end
		32'h0000067C: begin
				q			<=			16'h8067;
		end
		32'h0000067E: begin
				q			<=			16'h0000;
		end
		32'h00000680: begin
				q			<=			16'h0713;
		end
		32'h00000682: begin
				q			<=			16'h0010;
		end
		32'h00000684: begin
				q			<=			16'h8463;
		end
		32'h00000686: begin
				q			<=			16'h00E7;
		end
		32'h00000688: begin
				q			<=			16'h8067;
		end
		32'h0000068A: begin
				q			<=			16'h0000;
		end
		32'h0000068C: begin
				q			<=			16'h0713;
		end
		32'h0000068E: begin
				q			<=			16'h0000;
		end
		32'h00000690: begin
				q			<=			16'h15B7;
		end
		32'h00000692: begin
				q			<=			16'h0001;
		end
		32'h00000694: begin
				q			<=			16'h0637;
		end
		32'h00000696: begin
				q			<=			16'h4000;
		end
		32'h00000698: begin
				q			<=			16'h66B7;
		end
		32'h0000069A: begin
				q			<=			16'h0009;
		end
		32'h0000069C: begin
				q			<=			16'hA783;
		end
		32'h0000069E: begin
				q			<=			16'hF7C5;
		end
		32'h000006A0: begin
				q			<=			16'h07B3;
		end
		32'h000006A2: begin
				q			<=			16'h00F7;
		end
		32'h000006A4: begin
				q			<=			16'hE7B3;
		end
		32'h000006A6: begin
				q			<=			16'h00C7;
		end
		32'h000006A8: begin
				q			<=			16'hA023;
		end
		32'h000006AA: begin
				q			<=			16'h0007;
		end
		32'h000006AC: begin
				q			<=			16'h0713;
		end
		32'h000006AE: begin
				q			<=			16'h0047;
		end
		32'h000006B0: begin
				q			<=			16'h16E3;
		end
		32'h000006B2: begin
				q			<=			16'hFED7;
		end
		32'h000006B4: begin
				q			<=			16'hF06F;
		end
		32'h000006B6: begin
				q			<=			16'hFD5F;
		end
		32'h000006B8: begin
				q			<=			16'h0000;
		end
		32'h000006BA: begin
				q			<=			16'h0000;
		end
		32'h000006BC: begin
				q			<=			16'h17B7;
		end
		32'h000006BE: begin
				q			<=			16'h0001;
		end
		32'h000006C0: begin
				q			<=			16'hA783;
		end
		32'h000006C2: begin
				q			<=			16'hF787;
		end
		32'h000006C4: begin
				q			<=			16'h9A63;
		end
		32'h000006C6: begin
				q			<=			16'h0207;
		end
		32'h000006C8: begin
				q			<=			16'h0713;
		end
		32'h000006CA: begin
				q			<=			16'h0000;
		end
		32'h000006CC: begin
				q			<=			16'h1537;
		end
		32'h000006CE: begin
				q			<=			16'h0001;
		end
		32'h000006D0: begin
				q			<=			16'h05B7;
		end
		32'h000006D2: begin
				q			<=			16'h4000;
		end
		32'h000006D4: begin
				q			<=			16'h0613;
		end
		32'h000006D6: begin
				q			<=			16'hFFF0;
		end
		32'h000006D8: begin
				q			<=			16'h66B7;
		end
		32'h000006DA: begin
				q			<=			16'h0009;
		end
		32'h000006DC: begin
				q			<=			16'h2783;
		end
		32'h000006DE: begin
				q			<=			16'hF805;
		end
		32'h000006E0: begin
				q			<=			16'h07B3;
		end
		32'h000006E2: begin
				q			<=			16'h00F7;
		end
		32'h000006E4: begin
				q			<=			16'hE7B3;
		end
		32'h000006E6: begin
				q			<=			16'h00B7;
		end
		32'h000006E8: begin
				q			<=			16'hA023;
		end
		32'h000006EA: begin
				q			<=			16'h00C7;
		end
		32'h000006EC: begin
				q			<=			16'h0713;
		end
		32'h000006EE: begin
				q			<=			16'h0047;
		end
		32'h000006F0: begin
				q			<=			16'h16E3;
		end
		32'h000006F2: begin
				q			<=			16'hFED7;
		end
		32'h000006F4: begin
				q			<=			16'h8067;
		end
		32'h000006F6: begin
				q			<=			16'h0000;
		end
		32'h000006F8: begin
				q			<=			16'h0713;
		end
		32'h000006FA: begin
				q			<=			16'h0010;
		end
		32'h000006FC: begin
				q			<=			16'h8463;
		end
		32'h000006FE: begin
				q			<=			16'h00E7;
		end
		32'h00000700: begin
				q			<=			16'h8067;
		end
		32'h00000702: begin
				q			<=			16'h0000;
		end
		32'h00000704: begin
				q			<=			16'h0713;
		end
		32'h00000706: begin
				q			<=			16'h0000;
		end
		32'h00000708: begin
				q			<=			16'h1537;
		end
		32'h0000070A: begin
				q			<=			16'h0001;
		end
		32'h0000070C: begin
				q			<=			16'h05B7;
		end
		32'h0000070E: begin
				q			<=			16'h4000;
		end
		32'h00000710: begin
				q			<=			16'h0613;
		end
		32'h00000712: begin
				q			<=			16'hFFF0;
		end
		32'h00000714: begin
				q			<=			16'h66B7;
		end
		32'h00000716: begin
				q			<=			16'h0009;
		end
		32'h00000718: begin
				q			<=			16'h2783;
		end
		32'h0000071A: begin
				q			<=			16'hF7C5;
		end
		32'h0000071C: begin
				q			<=			16'h07B3;
		end
		32'h0000071E: begin
				q			<=			16'h00F7;
		end
		32'h00000720: begin
				q			<=			16'hE7B3;
		end
		32'h00000722: begin
				q			<=			16'h00B7;
		end
		32'h00000724: begin
				q			<=			16'hA023;
		end
		32'h00000726: begin
				q			<=			16'h00C7;
		end
		32'h00000728: begin
				q			<=			16'h0713;
		end
		32'h0000072A: begin
				q			<=			16'h0047;
		end
		32'h0000072C: begin
				q			<=			16'h16E3;
		end
		32'h0000072E: begin
				q			<=			16'hFED7;
		end
		32'h00000730: begin
				q			<=			16'hF06F;
		end
		32'h00000732: begin
				q			<=			16'hFD1F;
		end
		32'h00000734: begin
				q			<=			16'h0000;
		end
		32'h00000736: begin
				q			<=			16'h0000;
		end
		32'h00000738: begin
				q			<=			16'h0113;
		end
		32'h0000073A: begin
				q			<=			16'hFF01;
		end
		32'h0000073C: begin
				q			<=			16'h2623;
		end
		32'h0000073E: begin
				q			<=			16'h0011;
		end
		32'h00000740: begin
				q			<=			16'h0593;
		end
		32'h00000742: begin
				q			<=			16'h0010;
		end
		32'h00000744: begin
				q			<=			16'h0537;
		end
		32'h00000746: begin
				q			<=			16'h0001;
		end
		32'h00000748: begin
				q			<=			16'h0513;
		end
		32'h0000074A: begin
				q			<=			16'hA6C5;
		end
		32'h0000074C: begin
				q			<=			16'h00EF;
		end
		32'h0000074E: begin
				q			<=			16'h44C0;
		end
		32'h00000750: begin
				q			<=			16'h0593;
		end
		32'h00000752: begin
				q			<=			16'h0010;
		end
		32'h00000754: begin
				q			<=			16'h0537;
		end
		32'h00000756: begin
				q			<=			16'h0001;
		end
		32'h00000758: begin
				q			<=			16'h0513;
		end
		32'h0000075A: begin
				q			<=			16'hA845;
		end
		32'h0000075C: begin
				q			<=			16'h00EF;
		end
		32'h0000075E: begin
				q			<=			16'h43C0;
		end
		32'h00000760: begin
				q			<=			16'h0593;
		end
		32'h00000762: begin
				q			<=			16'h0010;
		end
		32'h00000764: begin
				q			<=			16'h0537;
		end
		32'h00000766: begin
				q			<=			16'h0001;
		end
		32'h00000768: begin
				q			<=			16'h0513;
		end
		32'h0000076A: begin
				q			<=			16'hAA85;
		end
		32'h0000076C: begin
				q			<=			16'h00EF;
		end
		32'h0000076E: begin
				q			<=			16'h42C0;
		end
		32'h00000770: begin
				q			<=			16'h0593;
		end
		32'h00000772: begin
				q			<=			16'h0010;
		end
		32'h00000774: begin
				q			<=			16'h0537;
		end
		32'h00000776: begin
				q			<=			16'h0001;
		end
		32'h00000778: begin
				q			<=			16'h0513;
		end
		32'h0000077A: begin
				q			<=			16'hAC85;
		end
		32'h0000077C: begin
				q			<=			16'h00EF;
		end
		32'h0000077E: begin
				q			<=			16'h41C0;
		end
		32'h00000780: begin
				q			<=			16'h0593;
		end
		32'h00000782: begin
				q			<=			16'h0010;
		end
		32'h00000784: begin
				q			<=			16'h0537;
		end
		32'h00000786: begin
				q			<=			16'h0001;
		end
		32'h00000788: begin
				q			<=			16'h0513;
		end
		32'h0000078A: begin
				q			<=			16'hAE85;
		end
		32'h0000078C: begin
				q			<=			16'h00EF;
		end
		32'h0000078E: begin
				q			<=			16'h40C0;
		end
		32'h00000790: begin
				q			<=			16'h0593;
		end
		32'h00000792: begin
				q			<=			16'h0010;
		end
		32'h00000794: begin
				q			<=			16'h0537;
		end
		32'h00000796: begin
				q			<=			16'h0001;
		end
		32'h00000798: begin
				q			<=			16'h0513;
		end
		32'h0000079A: begin
				q			<=			16'hB145;
		end
		32'h0000079C: begin
				q			<=			16'h00EF;
		end
		32'h0000079E: begin
				q			<=			16'h3FC0;
		end
		32'h000007A0: begin
				q			<=			16'h0593;
		end
		32'h000007A2: begin
				q			<=			16'h0010;
		end
		32'h000007A4: begin
				q			<=			16'h0537;
		end
		32'h000007A6: begin
				q			<=			16'h0001;
		end
		32'h000007A8: begin
				q			<=			16'h0513;
		end
		32'h000007AA: begin
				q			<=			16'hB405;
		end
		32'h000007AC: begin
				q			<=			16'h00EF;
		end
		32'h000007AE: begin
				q			<=			16'h3EC0;
		end
		32'h000007B0: begin
				q			<=			16'h0593;
		end
		32'h000007B2: begin
				q			<=			16'h0010;
		end
		32'h000007B4: begin
				q			<=			16'h0537;
		end
		32'h000007B6: begin
				q			<=			16'h0001;
		end
		32'h000007B8: begin
				q			<=			16'h0513;
		end
		32'h000007BA: begin
				q			<=			16'hB685;
		end
		32'h000007BC: begin
				q			<=			16'h00EF;
		end
		32'h000007BE: begin
				q			<=			16'h3DC0;
		end
		32'h000007C0: begin
				q			<=			16'h0593;
		end
		32'h000007C2: begin
				q			<=			16'h0010;
		end
		32'h000007C4: begin
				q			<=			16'h0537;
		end
		32'h000007C6: begin
				q			<=			16'h0001;
		end
		32'h000007C8: begin
				q			<=			16'h0513;
		end
		32'h000007CA: begin
				q			<=			16'hB8C5;
		end
		32'h000007CC: begin
				q			<=			16'h00EF;
		end
		32'h000007CE: begin
				q			<=			16'h3CC0;
		end
		32'h000007D0: begin
				q			<=			16'h2083;
		end
		32'h000007D2: begin
				q			<=			16'h00C1;
		end
		32'h000007D4: begin
				q			<=			16'h0113;
		end
		32'h000007D6: begin
				q			<=			16'h0101;
		end
		32'h000007D8: begin
				q			<=			16'h8067;
		end
		32'h000007DA: begin
				q			<=			16'h0000;
		end
		32'h000007DC: begin
				q			<=			16'h0000;
		end
		32'h000007DE: begin
				q			<=			16'h0000;
		end
		32'h000007E0: begin
				q			<=			16'h07B7;
		end
		32'h000007E2: begin
				q			<=			16'h8000;
		end
		32'h000007E4: begin
				q			<=			16'hA783;
		end
		32'h000007E6: begin
				q			<=			16'h0247;
		end
		32'h000007E8: begin
				q			<=			16'hF693;
		end
		32'h000007EA: begin
				q			<=			16'h0017;
		end
		32'h000007EC: begin
				q			<=			16'hE713;
		end
		32'h000007EE: begin
				q			<=			16'h0017;
		end
		32'h000007F0: begin
				q			<=			16'h9863;
		end
		32'h000007F2: begin
				q			<=			16'h0006;
		end
		32'h000007F4: begin
				q			<=			16'h07B7;
		end
		32'h000007F6: begin
				q			<=			16'h8000;
		end
		32'h000007F8: begin
				q			<=			16'hA223;
		end
		32'h000007FA: begin
				q			<=			16'h02E7;
		end
		32'h000007FC: begin
				q			<=			16'h8067;
		end
		32'h000007FE: begin
				q			<=			16'h0000;
		end
		32'h00000800: begin
				q			<=			16'hF713;
		end
		32'h00000802: begin
				q			<=			16'hFFE7;
		end
		32'h00000804: begin
				q			<=			16'hF06F;
		end
		32'h00000806: begin
				q			<=			16'hFF1F;
		end
		32'h00000808: begin
				q			<=			16'h0000;
		end
		32'h0000080A: begin
				q			<=			16'h0000;
		end
		32'h0000080C: begin
				q			<=			16'h0737;
		end
		32'h0000080E: begin
				q			<=			16'h8000;
		end
		32'h00000810: begin
				q			<=			16'h2783;
		end
		32'h00000812: begin
				q			<=			16'h0247;
		end
		32'h00000814: begin
				q			<=			16'hE793;
		end
		32'h00000816: begin
				q			<=			16'h0017;
		end
		32'h00000818: begin
				q			<=			16'h2223;
		end
		32'h0000081A: begin
				q			<=			16'h02F7;
		end
		32'h0000081C: begin
				q			<=			16'h8067;
		end
		32'h0000081E: begin
				q			<=			16'h0000;
		end
		32'h00000820: begin
				q			<=			16'h0000;
		end
		32'h00000822: begin
				q			<=			16'h0000;
		end
		32'h00000824: begin
				q			<=			16'h0737;
		end
		32'h00000826: begin
				q			<=			16'h8000;
		end
		32'h00000828: begin
				q			<=			16'h2783;
		end
		32'h0000082A: begin
				q			<=			16'h0247;
		end
		32'h0000082C: begin
				q			<=			16'hF793;
		end
		32'h0000082E: begin
				q			<=			16'hFFE7;
		end
		32'h00000830: begin
				q			<=			16'h2223;
		end
		32'h00000832: begin
				q			<=			16'h02F7;
		end
		32'h00000834: begin
				q			<=			16'h8067;
		end
		32'h00000836: begin
				q			<=			16'h0000;
		end
		32'h00000838: begin
				q			<=			16'h0000;
		end
		32'h0000083A: begin
				q			<=			16'h0000;
		end
		32'h0000083C: begin
				q			<=			16'h0113;
		end
		32'h0000083E: begin
				q			<=			16'hFF01;
		end
		32'h00000840: begin
				q			<=			16'h2623;
		end
		32'h00000842: begin
				q			<=			16'h0011;
		end
		32'h00000844: begin
				q			<=			16'h2423;
		end
		32'h00000846: begin
				q			<=			16'h0081;
		end
		32'h00000848: begin
				q			<=			16'h2223;
		end
		32'h0000084A: begin
				q			<=			16'h0091;
		end
		32'h0000084C: begin
				q			<=			16'h0613;
		end
		32'h0000084E: begin
				q			<=			16'h0040;
		end
		32'h00000850: begin
				q			<=			16'h05B7;
		end
		32'h00000852: begin
				q			<=			16'h0001;
		end
		32'h00000854: begin
				q			<=			16'h8593;
		end
		32'h00000856: begin
				q			<=			16'hBB05;
		end
		32'h00000858: begin
				q			<=			16'h1537;
		end
		32'h0000085A: begin
				q			<=			16'h0001;
		end
		32'h0000085C: begin
				q			<=			16'h0513;
		end
		32'h0000085E: begin
				q			<=			16'hC1C5;
		end
		32'h00000860: begin
				q			<=			16'h20EF;
		end
		32'h00000862: begin
				q			<=			16'h5EC0;
		end
		32'h00000864: begin
				q			<=			16'h0A63;
		end
		32'h00000866: begin
				q			<=			16'h0A05;
		end
		32'h00000868: begin
				q			<=			16'h0613;
		end
		32'h0000086A: begin
				q			<=			16'h0030;
		end
		32'h0000086C: begin
				q			<=			16'h05B7;
		end
		32'h0000086E: begin
				q			<=			16'h0001;
		end
		32'h00000870: begin
				q			<=			16'h8593;
		end
		32'h00000872: begin
				q			<=			16'hBB85;
		end
		32'h00000874: begin
				q			<=			16'h1537;
		end
		32'h00000876: begin
				q			<=			16'h0001;
		end
		32'h00000878: begin
				q			<=			16'h0513;
		end
		32'h0000087A: begin
				q			<=			16'hC1C5;
		end
		32'h0000087C: begin
				q			<=			16'h20EF;
		end
		32'h0000087E: begin
				q			<=			16'h5D00;
		end
		32'h00000880: begin
				q			<=			16'h0863;
		end
		32'h00000882: begin
				q			<=			16'h0A05;
		end
		32'h00000884: begin
				q			<=			16'h0613;
		end
		32'h00000886: begin
				q			<=			16'h0030;
		end
		32'h00000888: begin
				q			<=			16'h05B7;
		end
		32'h0000088A: begin
				q			<=			16'h0001;
		end
		32'h0000088C: begin
				q			<=			16'h8593;
		end
		32'h0000088E: begin
				q			<=			16'hBBC5;
		end
		32'h00000890: begin
				q			<=			16'h1537;
		end
		32'h00000892: begin
				q			<=			16'h0001;
		end
		32'h00000894: begin
				q			<=			16'h0513;
		end
		32'h00000896: begin
				q			<=			16'hC1C5;
		end
		32'h00000898: begin
				q			<=			16'h20EF;
		end
		32'h0000089A: begin
				q			<=			16'h5B40;
		end
		32'h0000089C: begin
				q			<=			16'h0E63;
		end
		32'h0000089E: begin
				q			<=			16'h0805;
		end
		32'h000008A0: begin
				q			<=			16'h0613;
		end
		32'h000008A2: begin
				q			<=			16'h0030;
		end
		32'h000008A4: begin
				q			<=			16'h05B7;
		end
		32'h000008A6: begin
				q			<=			16'h0001;
		end
		32'h000008A8: begin
				q			<=			16'h8593;
		end
		32'h000008AA: begin
				q			<=			16'hBC05;
		end
		32'h000008AC: begin
				q			<=			16'h1537;
		end
		32'h000008AE: begin
				q			<=			16'h0001;
		end
		32'h000008B0: begin
				q			<=			16'h0513;
		end
		32'h000008B2: begin
				q			<=			16'hC1C5;
		end
		32'h000008B4: begin
				q			<=			16'h20EF;
		end
		32'h000008B6: begin
				q			<=			16'h5980;
		end
		32'h000008B8: begin
				q			<=			16'h1E63;
		end
		32'h000008BA: begin
				q			<=			16'h0805;
		end
		32'h000008BC: begin
				q			<=			16'h14B7;
		end
		32'h000008BE: begin
				q			<=			16'h0001;
		end
		32'h000008C0: begin
				q			<=			16'h8513;
		end
		32'h000008C2: begin
				q			<=			16'hC1F4;
		end
		32'h000008C4: begin
				q			<=			16'h20EF;
		end
		32'h000008C6: begin
				q			<=			16'h5680;
		end
		32'h000008C8: begin
				q			<=			16'h0613;
		end
		32'h000008CA: begin
				q			<=			16'h0005;
		end
		32'h000008CC: begin
				q			<=			16'h1437;
		end
		32'h000008CE: begin
				q			<=			16'h0001;
		end
		32'h000008D0: begin
				q			<=			16'h0413;
		end
		32'h000008D2: begin
				q			<=			16'hF8C4;
		end
		32'h000008D4: begin
				q			<=			16'h2023;
		end
		32'h000008D6: begin
				q			<=			16'h00A4;
		end
		32'h000008D8: begin
				q			<=			16'h8593;
		end
		32'h000008DA: begin
				q			<=			16'hC1F4;
		end
		32'h000008DC: begin
				q			<=			16'h14B7;
		end
		32'h000008DE: begin
				q			<=			16'h0001;
		end
		32'h000008E0: begin
				q			<=			16'h8513;
		end
		32'h000008E2: begin
				q			<=			16'hB1C4;
		end
		32'h000008E4: begin
				q			<=			16'h20EF;
		end
		32'h000008E6: begin
				q			<=			16'h5A80;
		end
		32'h000008E8: begin
				q			<=			16'h2783;
		end
		32'h000008EA: begin
				q			<=			16'h0004;
		end
		32'h000008EC: begin
				q			<=			16'h8713;
		end
		32'h000008EE: begin
				q			<=			16'hB1C4;
		end
		32'h000008F0: begin
				q			<=			16'h87B3;
		end
		32'h000008F2: begin
				q			<=			16'h00E7;
		end
		32'h000008F4: begin
				q			<=			16'h8023;
		end
		32'h000008F6: begin
				q			<=			16'h0007;
		end
		32'h000008F8: begin
				q			<=			16'h8513;
		end
		32'h000008FA: begin
				q			<=			16'hB1C4;
		end
		32'h000008FC: begin
				q			<=			16'h10EF;
		end
		32'h000008FE: begin
				q			<=			16'h1700;
		end
		32'h00000900: begin
				q			<=			16'h1063;
		end
		32'h00000902: begin
				q			<=			16'h0405;
		end
		32'h00000904: begin
				q			<=			16'h0593;
		end
		32'h00000906: begin
				q			<=			16'h0010;
		end
		32'h00000908: begin
				q			<=			16'h0537;
		end
		32'h0000090A: begin
				q			<=			16'h0001;
		end
		32'h0000090C: begin
				q			<=			16'h0513;
		end
		32'h0000090E: begin
				q			<=			16'hBC45;
		end
		32'h00000910: begin
				q			<=			16'h00EF;
		end
		32'h00000912: begin
				q			<=			16'h2880;
		end
		32'h00000914: begin
				q			<=			16'h006F;
		end
		32'h00000916: begin
				q			<=			16'h0080;
		end
		32'h00000918: begin
				q			<=			16'hF0EF;
		end
		32'h0000091A: begin
				q			<=			16'hE21F;
		end
		32'h0000091C: begin
				q			<=			16'h2083;
		end
		32'h0000091E: begin
				q			<=			16'h00C1;
		end
		32'h00000920: begin
				q			<=			16'h2403;
		end
		32'h00000922: begin
				q			<=			16'h0081;
		end
		32'h00000924: begin
				q			<=			16'h2483;
		end
		32'h00000926: begin
				q			<=			16'h0041;
		end
		32'h00000928: begin
				q			<=			16'h0113;
		end
		32'h0000092A: begin
				q			<=			16'h0101;
		end
		32'h0000092C: begin
				q			<=			16'h8067;
		end
		32'h0000092E: begin
				q			<=			16'h0000;
		end
		32'h00000930: begin
				q			<=			16'h00EF;
		end
		32'h00000932: begin
				q			<=			16'h39C0;
		end
		32'h00000934: begin
				q			<=			16'hF06F;
		end
		32'h00000936: begin
				q			<=			16'hFE9F;
		end
		32'h00000938: begin
				q			<=			16'h10EF;
		end
		32'h0000093A: begin
				q			<=			16'h1C80;
		end
		32'h0000093C: begin
				q			<=			16'hF06F;
		end
		32'h0000093E: begin
				q			<=			16'hFE1F;
		end
		32'h00000940: begin
				q			<=			16'h0593;
		end
		32'h00000942: begin
				q			<=			16'h0010;
		end
		32'h00000944: begin
				q			<=			16'h0537;
		end
		32'h00000946: begin
				q			<=			16'h0001;
		end
		32'h00000948: begin
				q			<=			16'h0513;
		end
		32'h0000094A: begin
				q			<=			16'hBDC5;
		end
		32'h0000094C: begin
				q			<=			16'h00EF;
		end
		32'h0000094E: begin
				q			<=			16'h24C0;
		end
		32'h00000950: begin
				q			<=			16'hF06F;
		end
		32'h00000952: begin
				q			<=			16'hFCDF;
		end
		32'h00000954: begin
				q			<=			16'h0613;
		end
		32'h00000956: begin
				q			<=			16'h0080;
		end
		32'h00000958: begin
				q			<=			16'h05B7;
		end
		32'h0000095A: begin
				q			<=			16'h0001;
		end
		32'h0000095C: begin
				q			<=			16'h8593;
		end
		32'h0000095E: begin
				q			<=			16'hBF45;
		end
		32'h00000960: begin
				q			<=			16'h1537;
		end
		32'h00000962: begin
				q			<=			16'h0001;
		end
		32'h00000964: begin
				q			<=			16'h0513;
		end
		32'h00000966: begin
				q			<=			16'hC1C5;
		end
		32'h00000968: begin
				q			<=			16'h20EF;
		end
		32'h0000096A: begin
				q			<=			16'h4E40;
		end
		32'h0000096C: begin
				q			<=			16'h0063;
		end
		32'h0000096E: begin
				q			<=			16'h0A05;
		end
		32'h00000970: begin
				q			<=			16'h0613;
		end
		32'h00000972: begin
				q			<=			16'h0080;
		end
		32'h00000974: begin
				q			<=			16'h05B7;
		end
		32'h00000976: begin
				q			<=			16'h0001;
		end
		32'h00000978: begin
				q			<=			16'h8593;
		end
		32'h0000097A: begin
				q			<=			16'hC105;
		end
		32'h0000097C: begin
				q			<=			16'h1537;
		end
		32'h0000097E: begin
				q			<=			16'h0001;
		end
		32'h00000980: begin
				q			<=			16'h0513;
		end
		32'h00000982: begin
				q			<=			16'hC1C5;
		end
		32'h00000984: begin
				q			<=			16'h20EF;
		end
		32'h00000986: begin
				q			<=			16'h4C80;
		end
		32'h00000988: begin
				q			<=			16'h0E63;
		end
		32'h0000098A: begin
				q			<=			16'h0805;
		end
		32'h0000098C: begin
				q			<=			16'h0613;
		end
		32'h0000098E: begin
				q			<=			16'h0070;
		end
		32'h00000990: begin
				q			<=			16'h05B7;
		end
		32'h00000992: begin
				q			<=			16'h0001;
		end
		32'h00000994: begin
				q			<=			16'h8593;
		end
		32'h00000996: begin
				q			<=			16'hC2C5;
		end
		32'h00000998: begin
				q			<=			16'h1537;
		end
		32'h0000099A: begin
				q			<=			16'h0001;
		end
		32'h0000099C: begin
				q			<=			16'h0513;
		end
		32'h0000099E: begin
				q			<=			16'hC1C5;
		end
		32'h000009A0: begin
				q			<=			16'h20EF;
		end
		32'h000009A2: begin
				q			<=			16'h4AC0;
		end
		32'h000009A4: begin
				q			<=			16'h0C63;
		end
		32'h000009A6: begin
				q			<=			16'h0805;
		end
		32'h000009A8: begin
				q			<=			16'h0613;
		end
		32'h000009AA: begin
				q			<=			16'h0060;
		end
		32'h000009AC: begin
				q			<=			16'h05B7;
		end
		32'h000009AE: begin
				q			<=			16'h0001;
		end
		32'h000009B0: begin
				q			<=			16'h8593;
		end
		32'h000009B2: begin
				q			<=			16'hC445;
		end
		32'h000009B4: begin
				q			<=			16'h1537;
		end
		32'h000009B6: begin
				q			<=			16'h0001;
		end
		32'h000009B8: begin
				q			<=			16'h0513;
		end
		32'h000009BA: begin
				q			<=			16'hC1C5;
		end
		32'h000009BC: begin
				q			<=			16'h20EF;
		end
		32'h000009BE: begin
				q			<=			16'h4900;
		end
		32'h000009C0: begin
				q			<=			16'h0A63;
		end
		32'h000009C2: begin
				q			<=			16'h0805;
		end
		32'h000009C4: begin
				q			<=			16'h0613;
		end
		32'h000009C6: begin
				q			<=			16'h0070;
		end
		32'h000009C8: begin
				q			<=			16'h05B7;
		end
		32'h000009CA: begin
				q			<=			16'h0001;
		end
		32'h000009CC: begin
				q			<=			16'h8593;
		end
		32'h000009CE: begin
				q			<=			16'hC4C5;
		end
		32'h000009D0: begin
				q			<=			16'h1537;
		end
		32'h000009D2: begin
				q			<=			16'h0001;
		end
		32'h000009D4: begin
				q			<=			16'h0513;
		end
		32'h000009D6: begin
				q			<=			16'hC1C5;
		end
		32'h000009D8: begin
				q			<=			16'h20EF;
		end
		32'h000009DA: begin
				q			<=			16'h4740;
		end
		32'h000009DC: begin
				q			<=			16'h1463;
		end
		32'h000009DE: begin
				q			<=			16'h0A05;
		end
		32'h000009E0: begin
				q			<=			16'h17B7;
		end
		32'h000009E2: begin
				q			<=			16'h0001;
		end
		32'h000009E4: begin
				q			<=			16'hA783;
		end
		32'h000009E6: begin
				q			<=			16'hF787;
		end
		32'h000009E8: begin
				q			<=			16'h8263;
		end
		32'h000009EA: begin
				q			<=			16'h0807;
		end
		32'h000009EC: begin
				q			<=			16'h0713;
		end
		32'h000009EE: begin
				q			<=			16'h0010;
		end
		32'h000009F0: begin
				q			<=			16'h96E3;
		end
		32'h000009F2: begin
				q			<=			16'hF2E7;
		end
		32'h000009F4: begin
				q			<=			16'hF0EF;
		end
		32'h000009F6: begin
				q			<=			16'hBA1F;
		end
		32'h000009F8: begin
				q			<=			16'h0593;
		end
		32'h000009FA: begin
				q			<=			16'h0010;
		end
		32'h000009FC: begin
				q			<=			16'h0537;
		end
		32'h000009FE: begin
				q			<=			16'h0001;
		end
		32'h00000A00: begin
				q			<=			16'h0513;
		end
		32'h00000A02: begin
				q			<=			16'hC685;
		end
		32'h00000A04: begin
				q			<=			16'h00EF;
		end
		32'h00000A06: begin
				q			<=			16'h1940;
		end
		32'h00000A08: begin
				q			<=			16'hF06F;
		end
		32'h00000A0A: begin
				q			<=			16'hF15F;
		end
		32'h00000A0C: begin
				q			<=			16'hF0EF;
		end
		32'h00000A0E: begin
				q			<=			16'hC3DF;
		end
		32'h00000A10: begin
				q			<=			16'h0593;
		end
		32'h00000A12: begin
				q			<=			16'h0010;
		end
		32'h00000A14: begin
				q			<=			16'h0537;
		end
		32'h00000A16: begin
				q			<=			16'h0001;
		end
		32'h00000A18: begin
				q			<=			16'h0513;
		end
		32'h00000A1A: begin
				q			<=			16'hC005;
		end
		32'h00000A1C: begin
				q			<=			16'h00EF;
		end
		32'h00000A1E: begin
				q			<=			16'h17C0;
		end
		32'h00000A20: begin
				q			<=			16'hF06F;
		end
		32'h00000A22: begin
				q			<=			16'hEFDF;
		end
		32'h00000A24: begin
				q			<=			16'hF0EF;
		end
		32'h00000A26: begin
				q			<=			16'hC99F;
		end
		32'h00000A28: begin
				q			<=			16'h0593;
		end
		32'h00000A2A: begin
				q			<=			16'h0010;
		end
		32'h00000A2C: begin
				q			<=			16'h0537;
		end
		32'h00000A2E: begin
				q			<=			16'h0001;
		end
		32'h00000A30: begin
				q			<=			16'h0513;
		end
		32'h00000A32: begin
				q			<=			16'hC1C5;
		end
		32'h00000A34: begin
				q			<=			16'h00EF;
		end
		32'h00000A36: begin
				q			<=			16'h1640;
		end
		32'h00000A38: begin
				q			<=			16'hF06F;
		end
		32'h00000A3A: begin
				q			<=			16'hEE5F;
		end
		32'h00000A3C: begin
				q			<=			16'hF0EF;
		end
		32'h00000A3E: begin
				q			<=			16'hBA9F;
		end
		32'h00000A40: begin
				q			<=			16'h0593;
		end
		32'h00000A42: begin
				q			<=			16'h0010;
		end
		32'h00000A44: begin
				q			<=			16'h0537;
		end
		32'h00000A46: begin
				q			<=			16'h0001;
		end
		32'h00000A48: begin
				q			<=			16'h0513;
		end
		32'h00000A4A: begin
				q			<=			16'hC345;
		end
		32'h00000A4C: begin
				q			<=			16'h00EF;
		end
		32'h00000A4E: begin
				q			<=			16'h14C0;
		end
		32'h00000A50: begin
				q			<=			16'hF06F;
		end
		32'h00000A52: begin
				q			<=			16'hECDF;
		end
		32'h00000A54: begin
				q			<=			16'hF0EF;
		end
		32'h00000A56: begin
				q			<=			16'hB7DF;
		end
		32'h00000A58: begin
				q			<=			16'h0593;
		end
		32'h00000A5A: begin
				q			<=			16'h0010;
		end
		32'h00000A5C: begin
				q			<=			16'h0537;
		end
		32'h00000A5E: begin
				q			<=			16'h0001;
		end
		32'h00000A60: begin
				q			<=			16'h0513;
		end
		32'h00000A62: begin
				q			<=			16'hC345;
		end
		32'h00000A64: begin
				q			<=			16'h00EF;
		end
		32'h00000A66: begin
				q			<=			16'h1340;
		end
		32'h00000A68: begin
				q			<=			16'hF06F;
		end
		32'h00000A6A: begin
				q			<=			16'hEB5F;
		end
		32'h00000A6C: begin
				q			<=			16'hF0EF;
		end
		32'h00000A6E: begin
				q			<=			16'hB29F;
		end
		32'h00000A70: begin
				q			<=			16'h0593;
		end
		32'h00000A72: begin
				q			<=			16'h0010;
		end
		32'h00000A74: begin
				q			<=			16'h0537;
		end
		32'h00000A76: begin
				q			<=			16'h0001;
		end
		32'h00000A78: begin
				q			<=			16'h0513;
		end
		32'h00000A7A: begin
				q			<=			16'hC545;
		end
		32'h00000A7C: begin
				q			<=			16'h00EF;
		end
		32'h00000A7E: begin
				q			<=			16'h11C0;
		end
		32'h00000A80: begin
				q			<=			16'hF06F;
		end
		32'h00000A82: begin
				q			<=			16'hE9DF;
		end
		32'h00000A84: begin
				q			<=			16'h0613;
		end
		32'h00000A86: begin
				q			<=			16'h0060;
		end
		32'h00000A88: begin
				q			<=			16'h05B7;
		end
		32'h00000A8A: begin
				q			<=			16'h0001;
		end
		32'h00000A8C: begin
				q			<=			16'h8593;
		end
		32'h00000A8E: begin
				q			<=			16'hC7C5;
		end
		32'h00000A90: begin
				q			<=			16'h1537;
		end
		32'h00000A92: begin
				q			<=			16'h0001;
		end
		32'h00000A94: begin
				q			<=			16'h0513;
		end
		32'h00000A96: begin
				q			<=			16'hC1C5;
		end
		32'h00000A98: begin
				q			<=			16'h20EF;
		end
		32'h00000A9A: begin
				q			<=			16'h3B40;
		end
		32'h00000A9C: begin
				q			<=			16'h10E3;
		end
		32'h00000A9E: begin
				q			<=			16'hE805;
		end
		32'h00000AA0: begin
				q			<=			16'h07B7;
		end
		32'h00000AA2: begin
				q			<=			16'h8000;
		end
		32'h00000AA4: begin
				q			<=			16'hA403;
		end
		32'h00000AA6: begin
				q			<=			16'h0107;
		end
		32'h00000AA8: begin
				q			<=			16'h0593;
		end
		32'h00000AAA: begin
				q			<=			16'h0000;
		end
		32'h00000AAC: begin
				q			<=			16'h0537;
		end
		32'h00000AAE: begin
				q			<=			16'h0001;
		end
		32'h00000AB0: begin
				q			<=			16'h0513;
		end
		32'h00000AB2: begin
				q			<=			16'hC845;
		end
		32'h00000AB4: begin
				q			<=			16'h00EF;
		end
		32'h00000AB6: begin
				q			<=			16'h0E40;
		end
		32'h00000AB8: begin
				q			<=			16'h0513;
		end
		32'h00000ABA: begin
				q			<=			16'h0004;
		end
		32'h00000ABC: begin
				q			<=			16'h00EF;
		end
		32'h00000ABE: begin
				q			<=			16'h2880;
		end
		32'h00000AC0: begin
				q			<=			16'h0593;
		end
		32'h00000AC2: begin
				q			<=			16'h0010;
		end
		32'h00000AC4: begin
				q			<=			16'h0537;
		end
		32'h00000AC6: begin
				q			<=			16'h0001;
		end
		32'h00000AC8: begin
				q			<=			16'h0513;
		end
		32'h00000ACA: begin
				q			<=			16'hC8C5;
		end
		32'h00000ACC: begin
				q			<=			16'h00EF;
		end
		32'h00000ACE: begin
				q			<=			16'h0CC0;
		end
		32'h00000AD0: begin
				q			<=			16'hF06F;
		end
		32'h00000AD2: begin
				q			<=			16'hE4DF;
		end
		32'h00000AD4: begin
				q			<=			16'h0000;
		end
		32'h00000AD6: begin
				q			<=			16'h0000;
		end
		32'h00000AD8: begin
				q			<=			16'h0113;
		end
		32'h00000ADA: begin
				q			<=			16'hFF01;
		end
		32'h00000ADC: begin
				q			<=			16'h2623;
		end
		32'h00000ADE: begin
				q			<=			16'h0011;
		end
		32'h00000AE0: begin
				q			<=			16'h2423;
		end
		32'h00000AE2: begin
				q			<=			16'h0081;
		end
		32'h00000AE4: begin
				q			<=			16'h0793;
		end
		32'h00000AE6: begin
				q			<=			16'h0FF0;
		end
		32'h00000AE8: begin
				q			<=			16'h0663;
		end
		32'h00000AEA: begin
				q			<=			16'h06F5;
		end
		32'h00000AEC: begin
				q			<=			16'h0413;
		end
		32'h00000AEE: begin
				q			<=			16'h0005;
		end
		32'h00000AF0: begin
				q			<=			16'h0793;
		end
		32'h00000AF2: begin
				q			<=			16'hFEF5;
		end
		32'h00000AF4: begin
				q			<=			16'hF793;
		end
		32'h00000AF6: begin
				q			<=			16'h0FF7;
		end
		32'h00000AF8: begin
				q			<=			16'h0713;
		end
		32'h00000AFA: begin
				q			<=			16'h0030;
		end
		32'h00000AFC: begin
				q			<=			16'h7E63;
		end
		32'h00000AFE: begin
				q			<=			16'h04F7;
		end
		32'h00000B00: begin
				q			<=			16'h0793;
		end
		32'h00000B02: begin
				q			<=			16'h00A0;
		end
		32'h00000B04: begin
				q			<=			16'h1263;
		end
		32'h00000B06: begin
				q			<=			16'h06F5;
		end
		32'h00000B08: begin
				q			<=			16'h17B7;
		end
		32'h00000B0A: begin
				q			<=			16'h0001;
		end
		32'h00000B0C: begin
				q			<=			16'hA783;
		end
		32'h00000B0E: begin
				q			<=			16'hF887;
		end
		32'h00000B10: begin
				q			<=			16'h1737;
		end
		32'h00000B12: begin
				q			<=			16'h0001;
		end
		32'h00000B14: begin
				q			<=			16'h0713;
		end
		32'h00000B16: begin
				q			<=			16'hC1C7;
		end
		32'h00000B18: begin
				q			<=			16'h8733;
		end
		32'h00000B1A: begin
				q			<=			16'h00E7;
		end
		32'h00000B1C: begin
				q			<=			16'h0023;
		end
		32'h00000B1E: begin
				q			<=			16'h0007;
		end
		32'h00000B20: begin
				q			<=			16'h0713;
		end
		32'h00000B22: begin
				q			<=			16'h0500;
		end
		32'h00000B24: begin
				q			<=			16'hF7B3;
		end
		32'h00000B26: begin
				q			<=			16'h02E7;
		end
		32'h00000B28: begin
				q			<=			16'h8793;
		end
		32'h00000B2A: begin
				q			<=			16'h0017;
		end
		32'h00000B2C: begin
				q			<=			16'h6C63;
		end
		32'h00000B2E: begin
				q			<=			16'h00F7;
		end
		32'h00000B30: begin
				q			<=			16'h06B7;
		end
		32'h00000B32: begin
				q			<=			16'h8000;
		end
		32'h00000B34: begin
				q			<=			16'h0713;
		end
		32'h00000B36: begin
				q			<=			16'h0510;
		end
		32'h00000B38: begin
				q			<=			16'hA023;
		end
		32'h00000B3A: begin
				q			<=			16'h0006;
		end
		32'h00000B3C: begin
				q			<=			16'h8793;
		end
		32'h00000B3E: begin
				q			<=			16'h0017;
		end
		32'h00000B40: begin
				q			<=			16'h9CE3;
		end
		32'h00000B42: begin
				q			<=			16'hFEE7;
		end
		32'h00000B44: begin
				q			<=			16'hF0EF;
		end
		32'h00000B46: begin
				q			<=			16'hCF9F;
		end
		32'h00000B48: begin
				q			<=			16'h17B7;
		end
		32'h00000B4A: begin
				q			<=			16'h0001;
		end
		32'h00000B4C: begin
				q			<=			16'hA423;
		end
		32'h00000B4E: begin
				q			<=			16'hF807;
		end
		32'h00000B50: begin
				q			<=			16'h006F;
		end
		32'h00000B52: begin
				q			<=			16'h0080;
		end
		32'h00000B54: begin
				q			<=			16'hF0EF;
		end
		32'h00000B56: begin
				q			<=			16'hC8DF;
		end
		32'h00000B58: begin
				q			<=			16'h2083;
		end
		32'h00000B5A: begin
				q			<=			16'h00C1;
		end
		32'h00000B5C: begin
				q			<=			16'h2403;
		end
		32'h00000B5E: begin
				q			<=			16'h0081;
		end
		32'h00000B60: begin
				q			<=			16'h0113;
		end
		32'h00000B62: begin
				q			<=			16'h0101;
		end
		32'h00000B64: begin
				q			<=			16'h8067;
		end
		32'h00000B66: begin
				q			<=			16'h0000;
		end
		32'h00000B68: begin
				q			<=			16'h00EF;
		end
		32'h00000B6A: begin
				q			<=			16'h1400;
		end
		32'h00000B6C: begin
				q			<=			16'h1737;
		end
		32'h00000B6E: begin
				q			<=			16'h0001;
		end
		32'h00000B70: begin
				q			<=			16'h0713;
		end
		32'h00000B72: begin
				q			<=			16'hF887;
		end
		32'h00000B74: begin
				q			<=			16'h2683;
		end
		32'h00000B76: begin
				q			<=			16'h0007;
		end
		32'h00000B78: begin
				q			<=			16'h17B7;
		end
		32'h00000B7A: begin
				q			<=			16'h0001;
		end
		32'h00000B7C: begin
				q			<=			16'h8793;
		end
		32'h00000B7E: begin
				q			<=			16'hC1C7;
		end
		32'h00000B80: begin
				q			<=			16'h87B3;
		end
		32'h00000B82: begin
				q			<=			16'h00F6;
		end
		32'h00000B84: begin
				q			<=			16'h8023;
		end
		32'h00000B86: begin
				q			<=			16'h0087;
		end
		32'h00000B88: begin
				q			<=			16'h8693;
		end
		32'h00000B8A: begin
				q			<=			16'h0016;
		end
		32'h00000B8C: begin
				q			<=			16'h2023;
		end
		32'h00000B8E: begin
				q			<=			16'h00D7;
		end
		32'h00000B90: begin
				q			<=			16'hF06F;
		end
		32'h00000B92: begin
				q			<=			16'hFC9F;
		end
		32'h00000B94: begin
				q			<=			16'h0000;
		end
		32'h00000B96: begin
				q			<=			16'h0000;
		end
		32'h00000B98: begin
				q			<=			16'h0113;
		end
		32'h00000B9A: begin
				q			<=			16'hFF01;
		end
		32'h00000B9C: begin
				q			<=			16'h2623;
		end
		32'h00000B9E: begin
				q			<=			16'h0011;
		end
		32'h00000BA0: begin
				q			<=			16'h2423;
		end
		32'h00000BA2: begin
				q			<=			16'h0081;
		end
		32'h00000BA4: begin
				q			<=			16'h2223;
		end
		32'h00000BA6: begin
				q			<=			16'h0091;
		end
		32'h00000BA8: begin
				q			<=			16'h0413;
		end
		32'h00000BAA: begin
				q			<=			16'h0005;
		end
		32'h00000BAC: begin
				q			<=			16'h8493;
		end
		32'h00000BAE: begin
				q			<=			16'h0005;
		end
		32'h00000BB0: begin
				q			<=			16'h20EF;
		end
		32'h00000BB2: begin
				q			<=			16'h27C0;
		end
		32'h00000BB4: begin
				q			<=			16'h0713;
		end
		32'h00000BB6: begin
				q			<=			16'h0004;
		end
		32'h00000BB8: begin
				q			<=			16'h0693;
		end
		32'h00000BBA: begin
				q			<=			16'h0000;
		end
		32'h00000BBC: begin
				q			<=			16'h0837;
		end
		32'h00000BBE: begin
				q			<=			16'h8000;
		end
		32'h00000BC0: begin
				q			<=			16'h15B7;
		end
		32'h00000BC2: begin
				q			<=			16'h0001;
		end
		32'h00000BC4: begin
				q			<=			16'h4783;
		end
		32'h00000BC6: begin
				q			<=			16'h0007;
		end
		32'h00000BC8: begin
				q			<=			16'h2023;
		end
		32'h00000BCA: begin
				q			<=			16'h00F8;
		end
		32'h00000BCC: begin
				q			<=			16'h8613;
		end
		32'h00000BCE: begin
				q			<=			16'hF905;
		end
		32'h00000BD0: begin
				q			<=			16'h2783;
		end
		32'h00000BD2: begin
				q			<=			16'h0006;
		end
		32'h00000BD4: begin
				q			<=			16'h8793;
		end
		32'h00000BD6: begin
				q			<=			16'h0017;
		end
		32'h00000BD8: begin
				q			<=			16'h2023;
		end
		32'h00000BDA: begin
				q			<=			16'h00F6;
		end
		32'h00000BDC: begin
				q			<=			16'h8693;
		end
		32'h00000BDE: begin
				q			<=			16'h0016;
		end
		32'h00000BE0: begin
				q			<=			16'h0713;
		end
		32'h00000BE2: begin
				q			<=			16'h0017;
		end
		32'h00000BE4: begin
				q			<=			16'h70E3;
		end
		32'h00000BE6: begin
				q			<=			16'hFED5;
		end
		32'h00000BE8: begin
				q			<=			16'h8063;
		end
		32'h00000BEA: begin
				q			<=			16'h0404;
		end
		32'h00000BEC: begin
				q			<=			16'h0793;
		end
		32'h00000BEE: begin
				q			<=			16'h0500;
		end
		32'h00000BF0: begin
				q			<=			16'h7533;
		end
		32'h00000BF2: begin
				q			<=			16'h02F5;
		end
		32'h00000BF4: begin
				q			<=			16'h0513;
		end
		32'h00000BF6: begin
				q			<=			16'h0015;
		end
		32'h00000BF8: begin
				q			<=			16'h0793;
		end
		32'h00000BFA: begin
				q			<=			16'h04F0;
		end
		32'h00000BFC: begin
				q			<=			16'hE663;
		end
		32'h00000BFE: begin
				q			<=			16'h02A7;
		end
		32'h00000C00: begin
				q			<=			16'h05B7;
		end
		32'h00000C02: begin
				q			<=			16'h8000;
		end
		32'h00000C04: begin
				q			<=			16'h1637;
		end
		32'h00000C06: begin
				q			<=			16'h0001;
		end
		32'h00000C08: begin
				q			<=			16'h0693;
		end
		32'h00000C0A: begin
				q			<=			16'h0500;
		end
		32'h00000C0C: begin
				q			<=			16'hA023;
		end
		32'h00000C0E: begin
				q			<=			16'h0005;
		end
		32'h00000C10: begin
				q			<=			16'h0713;
		end
		32'h00000C12: begin
				q			<=			16'hF906;
		end
		32'h00000C14: begin
				q			<=			16'h2783;
		end
		32'h00000C16: begin
				q			<=			16'h0007;
		end
		32'h00000C18: begin
				q			<=			16'h8793;
		end
		32'h00000C1A: begin
				q			<=			16'h0017;
		end
		32'h00000C1C: begin
				q			<=			16'h2023;
		end
		32'h00000C1E: begin
				q			<=			16'h00F7;
		end
		32'h00000C20: begin
				q			<=			16'h0513;
		end
		32'h00000C22: begin
				q			<=			16'h0015;
		end
		32'h00000C24: begin
				q			<=			16'h14E3;
		end
		32'h00000C26: begin
				q			<=			16'hFED5;
		end
		32'h00000C28: begin
				q			<=			16'h2083;
		end
		32'h00000C2A: begin
				q			<=			16'h00C1;
		end
		32'h00000C2C: begin
				q			<=			16'h2403;
		end
		32'h00000C2E: begin
				q			<=			16'h0081;
		end
		32'h00000C30: begin
				q			<=			16'h2483;
		end
		32'h00000C32: begin
				q			<=			16'h0041;
		end
		32'h00000C34: begin
				q			<=			16'h0113;
		end
		32'h00000C36: begin
				q			<=			16'h0101;
		end
		32'h00000C38: begin
				q			<=			16'h8067;
		end
		32'h00000C3A: begin
				q			<=			16'h0000;
		end
		32'h00000C3C: begin
				q			<=			16'h0000;
		end
		32'h00000C3E: begin
				q			<=			16'h0000;
		end
		32'h00000C40: begin
				q			<=			16'h0113;
		end
		32'h00000C42: begin
				q			<=			16'hDF01;
		end
		32'h00000C44: begin
				q			<=			16'h2623;
		end
		32'h00000C46: begin
				q			<=			16'h2011;
		end
		32'h00000C48: begin
				q			<=			16'h0713;
		end
		32'h00000C4A: begin
				q			<=			16'h0005;
		end
		32'h00000C4C: begin
				q			<=			16'h06B7;
		end
		32'h00000C4E: begin
				q			<=			16'h0001;
		end
		32'h00000C50: begin
				q			<=			16'h8693;
		end
		32'h00000C52: begin
				q			<=			16'hC906;
		end
		32'h00000C54: begin
				q			<=			16'h0637;
		end
		32'h00000C56: begin
				q			<=			16'h0001;
		end
		32'h00000C58: begin
				q			<=			16'h0613;
		end
		32'h00000C5A: begin
				q			<=			16'hC9C6;
		end
		32'h00000C5C: begin
				q			<=			16'h0593;
		end
		32'h00000C5E: begin
				q			<=			16'h2000;
		end
		32'h00000C60: begin
				q			<=			16'h0513;
		end
		32'h00000C62: begin
				q			<=			16'h0001;
		end
		32'h00000C64: begin
				q			<=			16'h2097;
		end
		32'h00000C66: begin
				q			<=			16'h0000;
		end
		32'h00000C68: begin
				q			<=			16'h80E7;
		end
		32'h00000C6A: begin
				q			<=			16'h1080;
		end
		32'h00000C6C: begin
				q			<=			16'h0593;
		end
		32'h00000C6E: begin
				q			<=			16'h0010;
		end
		32'h00000C70: begin
				q			<=			16'h0513;
		end
		32'h00000C72: begin
				q			<=			16'h0001;
		end
		32'h00000C74: begin
				q			<=			16'hF0EF;
		end
		32'h00000C76: begin
				q			<=			16'hF25F;
		end
		32'h00000C78: begin
				q			<=			16'h2083;
		end
		32'h00000C7A: begin
				q			<=			16'h20C1;
		end
		32'h00000C7C: begin
				q			<=			16'h0113;
		end
		32'h00000C7E: begin
				q			<=			16'h2101;
		end
		32'h00000C80: begin
				q			<=			16'h8067;
		end
		32'h00000C82: begin
				q			<=			16'h0000;
		end
		32'h00000C84: begin
				q			<=			16'h0000;
		end
		32'h00000C86: begin
				q			<=			16'h0000;
		end
		32'h00000C88: begin
				q			<=			16'h0113;
		end
		32'h00000C8A: begin
				q			<=			16'hFF01;
		end
		32'h00000C8C: begin
				q			<=			16'h2623;
		end
		32'h00000C8E: begin
				q			<=			16'h0011;
		end
		32'h00000C90: begin
				q			<=			16'h0593;
		end
		32'h00000C92: begin
				q			<=			16'h0010;
		end
		32'h00000C94: begin
				q			<=			16'hF0EF;
		end
		32'h00000C96: begin
				q			<=			16'hF05F;
		end
		32'h00000C98: begin
				q			<=			16'h2083;
		end
		32'h00000C9A: begin
				q			<=			16'h00C1;
		end
		32'h00000C9C: begin
				q			<=			16'h0113;
		end
		32'h00000C9E: begin
				q			<=			16'h0101;
		end
		32'h00000CA0: begin
				q			<=			16'h8067;
		end
		32'h00000CA2: begin
				q			<=			16'h0000;
		end
		32'h00000CA4: begin
				q			<=			16'h0000;
		end
		32'h00000CA6: begin
				q			<=			16'h0000;
		end
		32'h00000CA8: begin
				q			<=			16'h07B7;
		end
		32'h00000CAA: begin
				q			<=			16'h8000;
		end
		32'h00000CAC: begin
				q			<=			16'hA023;
		end
		32'h00000CAE: begin
				q			<=			16'h00A7;
		end
		32'h00000CB0: begin
				q			<=			16'h17B7;
		end
		32'h00000CB2: begin
				q			<=			16'h0001;
		end
		32'h00000CB4: begin
				q			<=			16'h8793;
		end
		32'h00000CB6: begin
				q			<=			16'hF907;
		end
		32'h00000CB8: begin
				q			<=			16'hA703;
		end
		32'h00000CBA: begin
				q			<=			16'h0007;
		end
		32'h00000CBC: begin
				q			<=			16'h0713;
		end
		32'h00000CBE: begin
				q			<=			16'h0017;
		end
		32'h00000CC0: begin
				q			<=			16'hA023;
		end
		32'h00000CC2: begin
				q			<=			16'h00E7;
		end
		32'h00000CC4: begin
				q			<=			16'h8067;
		end
		32'h00000CC6: begin
				q			<=			16'h0000;
		end
		32'h00000CC8: begin
				q			<=			16'h0000;
		end
		32'h00000CCA: begin
				q			<=			16'h0000;
		end
		32'h00000CCC: begin
				q			<=			16'h0737;
		end
		32'h00000CCE: begin
				q			<=			16'h8000;
		end
		32'h00000CD0: begin
				q			<=			16'h2783;
		end
		32'h00000CD2: begin
				q			<=			16'h0247;
		end
		32'h00000CD4: begin
				q			<=			16'hE793;
		end
		32'h00000CD6: begin
				q			<=			16'h0027;
		end
		32'h00000CD8: begin
				q			<=			16'h2223;
		end
		32'h00000CDA: begin
				q			<=			16'h02F7;
		end
		32'h00000CDC: begin
				q			<=			16'h17B7;
		end
		32'h00000CDE: begin
				q			<=			16'h0001;
		end
		32'h00000CE0: begin
				q			<=			16'hA823;
		end
		32'h00000CE2: begin
				q			<=			16'hF807;
		end
		32'h00000CE4: begin
				q			<=			16'h8067;
		end
		32'h00000CE6: begin
				q			<=			16'h0000;
		end
		32'h00000CE8: begin
				q			<=			16'h0000;
		end
		32'h00000CEA: begin
				q			<=			16'h0000;
		end
		32'h00000CEC: begin
				q			<=			16'h0737;
		end
		32'h00000CEE: begin
				q			<=			16'h8000;
		end
		32'h00000CF0: begin
				q			<=			16'h2783;
		end
		32'h00000CF2: begin
				q			<=			16'h0247;
		end
		32'h00000CF4: begin
				q			<=			16'hE793;
		end
		32'h00000CF6: begin
				q			<=			16'h0047;
		end
		32'h00000CF8: begin
				q			<=			16'h2223;
		end
		32'h00000CFA: begin
				q			<=			16'h02F7;
		end
		32'h00000CFC: begin
				q			<=			16'h17B7;
		end
		32'h00000CFE: begin
				q			<=			16'h0001;
		end
		32'h00000D00: begin
				q			<=			16'h8793;
		end
		32'h00000D02: begin
				q			<=			16'hF907;
		end
		32'h00000D04: begin
				q			<=			16'hA703;
		end
		32'h00000D06: begin
				q			<=			16'h0007;
		end
		32'h00000D08: begin
				q			<=			16'h0693;
		end
		32'h00000D0A: begin
				q			<=			16'h03C0;
		end
		32'h00000D0C: begin
				q			<=			16'h5733;
		end
		32'h00000D0E: begin
				q			<=			16'h02D7;
		end
		32'h00000D10: begin
				q			<=			16'hA023;
		end
		32'h00000D12: begin
				q			<=			16'h00E7;
		end
		32'h00000D14: begin
				q			<=			16'h8067;
		end
		32'h00000D16: begin
				q			<=			16'h0000;
		end
		32'h00000D18: begin
				q			<=			16'h0000;
		end
		32'h00000D1A: begin
				q			<=			16'h0000;
		end
		32'h00000D1C: begin
				q			<=			16'hD5B3;
		end
		32'h00000D1E: begin
				q			<=			16'h00A5;
		end
		32'h00000D20: begin
				q			<=			16'hF593;
		end
		32'h00000D22: begin
				q			<=			16'h0015;
		end
		32'h00000D24: begin
				q			<=			16'h9863;
		end
		32'h00000D26: begin
				q			<=			16'h0005;
		end
		32'h00000D28: begin
				q			<=			16'h1537;
		end
		32'h00000D2A: begin
				q			<=			16'h0001;
		end
		32'h00000D2C: begin
				q			<=			16'h0513;
		end
		32'h00000D2E: begin
				q			<=			16'h8E85;
		end
		32'h00000D30: begin
				q			<=			16'h8067;
		end
		32'h00000D32: begin
				q			<=			16'h0000;
		end
		32'h00000D34: begin
				q			<=			16'h1537;
		end
		32'h00000D36: begin
				q			<=			16'h0001;
		end
		32'h00000D38: begin
				q			<=			16'h0513;
		end
		32'h00000D3A: begin
				q			<=			16'h8E45;
		end
		32'h00000D3C: begin
				q			<=			16'h8067;
		end
		32'h00000D3E: begin
				q			<=			16'h0000;
		end
		32'h00000D40: begin
				q			<=			16'h0000;
		end
		32'h00000D42: begin
				q			<=			16'h0000;
		end
		32'h00000D44: begin
				q			<=			16'h0113;
		end
		32'h00000D46: begin
				q			<=			16'hFE01;
		end
		32'h00000D48: begin
				q			<=			16'h2E23;
		end
		32'h00000D4A: begin
				q			<=			16'h0011;
		end
		32'h00000D4C: begin
				q			<=			16'h2C23;
		end
		32'h00000D4E: begin
				q			<=			16'h0081;
		end
		32'h00000D50: begin
				q			<=			16'h0413;
		end
		32'h00000D52: begin
				q			<=			16'h0005;
		end
		32'h00000D54: begin
				q			<=			16'h4A63;
		end
		32'h00000D56: begin
				q			<=			16'h3005;
		end
		32'h00000D58: begin
				q			<=			16'h16B7;
		end
		32'h00000D5A: begin
				q			<=			16'h0001;
		end
		32'h00000D5C: begin
				q			<=			16'h8693;
		end
		32'h00000D5E: begin
				q			<=			16'h8E86;
		end
		32'h00000D60: begin
				q			<=			16'h1793;
		end
		32'h00000D62: begin
				q			<=			16'h0014;
		end
		32'h00000D64: begin
				q			<=			16'hC863;
		end
		32'h00000D66: begin
				q			<=			16'h3007;
		end
		32'h00000D68: begin
				q			<=			16'h1737;
		end
		32'h00000D6A: begin
				q			<=			16'h0001;
		end
		32'h00000D6C: begin
				q			<=			16'h0713;
		end
		32'h00000D6E: begin
				q			<=			16'h8E87;
		end
		32'h00000D70: begin
				q			<=			16'h1793;
		end
		32'h00000D72: begin
				q			<=			16'h0024;
		end
		32'h00000D74: begin
				q			<=			16'hC663;
		end
		32'h00000D76: begin
				q			<=			16'h3007;
		end
		32'h00000D78: begin
				q			<=			16'h17B7;
		end
		32'h00000D7A: begin
				q			<=			16'h0001;
		end
		32'h00000D7C: begin
				q			<=			16'h8793;
		end
		32'h00000D7E: begin
				q			<=			16'h8E87;
		end
		32'h00000D80: begin
				q			<=			16'h1613;
		end
		32'h00000D82: begin
				q			<=			16'h0034;
		end
		32'h00000D84: begin
				q			<=			16'h4463;
		end
		32'h00000D86: begin
				q			<=			16'h3006;
		end
		32'h00000D88: begin
				q			<=			16'h1837;
		end
		32'h00000D8A: begin
				q			<=			16'h0001;
		end
		32'h00000D8C: begin
				q			<=			16'h0813;
		end
		32'h00000D8E: begin
				q			<=			16'h8E88;
		end
		32'h00000D90: begin
				q			<=			16'h1613;
		end
		32'h00000D92: begin
				q			<=			16'h0044;
		end
		32'h00000D94: begin
				q			<=			16'h4263;
		end
		32'h00000D96: begin
				q			<=			16'h3006;
		end
		32'h00000D98: begin
				q			<=			16'h18B7;
		end
		32'h00000D9A: begin
				q			<=			16'h0001;
		end
		32'h00000D9C: begin
				q			<=			16'h8893;
		end
		32'h00000D9E: begin
				q			<=			16'h8E88;
		end
		32'h00000DA0: begin
				q			<=			16'h1613;
		end
		32'h00000DA2: begin
				q			<=			16'h0054;
		end
		32'h00000DA4: begin
				q			<=			16'h4063;
		end
		32'h00000DA6: begin
				q			<=			16'h3006;
		end
		32'h00000DA8: begin
				q			<=			16'h1637;
		end
		32'h00000DAA: begin
				q			<=			16'h0001;
		end
		32'h00000DAC: begin
				q			<=			16'h0613;
		end
		32'h00000DAE: begin
				q			<=			16'h8E86;
		end
		32'h00000DB0: begin
				q			<=			16'h1593;
		end
		32'h00000DB2: begin
				q			<=			16'h0064;
		end
		32'h00000DB4: begin
				q			<=			16'hCE63;
		end
		32'h00000DB6: begin
				q			<=			16'h2E05;
		end
		32'h00000DB8: begin
				q			<=			16'h15B7;
		end
		32'h00000DBA: begin
				q			<=			16'h0001;
		end
		32'h00000DBC: begin
				q			<=			16'h8593;
		end
		32'h00000DBE: begin
				q			<=			16'h8E85;
		end
		32'h00000DC0: begin
				q			<=			16'h1513;
		end
		32'h00000DC2: begin
				q			<=			16'h0074;
		end
		32'h00000DC4: begin
				q			<=			16'h4C63;
		end
		32'h00000DC6: begin
				q			<=			16'h2E05;
		end
		32'h00000DC8: begin
				q			<=			16'h1537;
		end
		32'h00000DCA: begin
				q			<=			16'h0001;
		end
		32'h00000DCC: begin
				q			<=			16'h0513;
		end
		32'h00000DCE: begin
				q			<=			16'h8E85;
		end
		32'h00000DD0: begin
				q			<=			16'h2423;
		end
		32'h00000DD2: begin
				q			<=			16'h00A1;
		end
		32'h00000DD4: begin
				q			<=			16'h2223;
		end
		32'h00000DD6: begin
				q			<=			16'h00B1;
		end
		32'h00000DD8: begin
				q			<=			16'h2023;
		end
		32'h00000DDA: begin
				q			<=			16'h00C1;
		end
		32'h00000DDC: begin
				q			<=			16'h0637;
		end
		32'h00000DDE: begin
				q			<=			16'h0001;
		end
		32'h00000DE0: begin
				q			<=			16'h0613;
		end
		32'h00000DE2: begin
				q			<=			16'hCA46;
		end
		32'h00000DE4: begin
				q			<=			16'h0593;
		end
		32'h00000DE6: begin
				q			<=			16'h1000;
		end
		32'h00000DE8: begin
				q			<=			16'h1537;
		end
		32'h00000DEA: begin
				q			<=			16'h0001;
		end
		32'h00000DEC: begin
				q			<=			16'h0513;
		end
		32'h00000DEE: begin
				q			<=			16'hD1C5;
		end
		32'h00000DF0: begin
				q			<=			16'h2097;
		end
		32'h00000DF2: begin
				q			<=			16'h0000;
		end
		32'h00000DF4: begin
				q			<=			16'h80E7;
		end
		32'h00000DF6: begin
				q			<=			16'hF7C0;
		end
		32'h00000DF8: begin
				q			<=			16'h1793;
		end
		32'h00000DFA: begin
				q			<=			16'h0084;
		end
		32'h00000DFC: begin
				q			<=			16'hC663;
		end
		32'h00000DFE: begin
				q			<=			16'h2C07;
		end
		32'h00000E00: begin
				q			<=			16'h1737;
		end
		32'h00000E02: begin
				q			<=			16'h0001;
		end
		32'h00000E04: begin
				q			<=			16'h0713;
		end
		32'h00000E06: begin
				q			<=			16'h8E87;
		end
		32'h00000E08: begin
				q			<=			16'h1793;
		end
		32'h00000E0A: begin
				q			<=			16'h0094;
		end
		32'h00000E0C: begin
				q			<=			16'hC463;
		end
		32'h00000E0E: begin
				q			<=			16'h2C07;
		end
		32'h00000E10: begin
				q			<=			16'h17B7;
		end
		32'h00000E12: begin
				q			<=			16'h0001;
		end
		32'h00000E14: begin
				q			<=			16'h8793;
		end
		32'h00000E16: begin
				q			<=			16'h8E87;
		end
		32'h00000E18: begin
				q			<=			16'h1693;
		end
		32'h00000E1A: begin
				q			<=			16'h00A4;
		end
		32'h00000E1C: begin
				q			<=			16'hC263;
		end
		32'h00000E1E: begin
				q			<=			16'h2C06;
		end
		32'h00000E20: begin
				q			<=			16'h1837;
		end
		32'h00000E22: begin
				q			<=			16'h0001;
		end
		32'h00000E24: begin
				q			<=			16'h0813;
		end
		32'h00000E26: begin
				q			<=			16'h8E88;
		end
		32'h00000E28: begin
				q			<=			16'h1693;
		end
		32'h00000E2A: begin
				q			<=			16'h00B4;
		end
		32'h00000E2C: begin
				q			<=			16'hC063;
		end
		32'h00000E2E: begin
				q			<=			16'h2C06;
		end
		32'h00000E30: begin
				q			<=			16'h18B7;
		end
		32'h00000E32: begin
				q			<=			16'h0001;
		end
		32'h00000E34: begin
				q			<=			16'h8893;
		end
		32'h00000E36: begin
				q			<=			16'h8E88;
		end
		32'h00000E38: begin
				q			<=			16'h1693;
		end
		32'h00000E3A: begin
				q			<=			16'h00C4;
		end
		32'h00000E3C: begin
				q			<=			16'hCE63;
		end
		32'h00000E3E: begin
				q			<=			16'h2A06;
		end
		32'h00000E40: begin
				q			<=			16'h16B7;
		end
		32'h00000E42: begin
				q			<=			16'h0001;
		end
		32'h00000E44: begin
				q			<=			16'h8693;
		end
		32'h00000E46: begin
				q			<=			16'h8E86;
		end
		32'h00000E48: begin
				q			<=			16'h1613;
		end
		32'h00000E4A: begin
				q			<=			16'h00D4;
		end
		32'h00000E4C: begin
				q			<=			16'h4C63;
		end
		32'h00000E4E: begin
				q			<=			16'h2A06;
		end
		32'h00000E50: begin
				q			<=			16'h1637;
		end
		32'h00000E52: begin
				q			<=			16'h0001;
		end
		32'h00000E54: begin
				q			<=			16'h0613;
		end
		32'h00000E56: begin
				q			<=			16'h8E86;
		end
		32'h00000E58: begin
				q			<=			16'h1593;
		end
		32'h00000E5A: begin
				q			<=			16'h00E4;
		end
		32'h00000E5C: begin
				q			<=			16'hCA63;
		end
		32'h00000E5E: begin
				q			<=			16'h2A05;
		end
		32'h00000E60: begin
				q			<=			16'h15B7;
		end
		32'h00000E62: begin
				q			<=			16'h0001;
		end
		32'h00000E64: begin
				q			<=			16'h8593;
		end
		32'h00000E66: begin
				q			<=			16'h8E85;
		end
		32'h00000E68: begin
				q			<=			16'h1513;
		end
		32'h00000E6A: begin
				q			<=			16'h00F4;
		end
		32'h00000E6C: begin
				q			<=			16'h4863;
		end
		32'h00000E6E: begin
				q			<=			16'h2A05;
		end
		32'h00000E70: begin
				q			<=			16'h1537;
		end
		32'h00000E72: begin
				q			<=			16'h0001;
		end
		32'h00000E74: begin
				q			<=			16'h0513;
		end
		32'h00000E76: begin
				q			<=			16'h8E85;
		end
		32'h00000E78: begin
				q			<=			16'h2623;
		end
		32'h00000E7A: begin
				q			<=			16'h00A1;
		end
		32'h00000E7C: begin
				q			<=			16'h2423;
		end
		32'h00000E7E: begin
				q			<=			16'h00B1;
		end
		32'h00000E80: begin
				q			<=			16'h2223;
		end
		32'h00000E82: begin
				q			<=			16'h00C1;
		end
		32'h00000E84: begin
				q			<=			16'h2023;
		end
		32'h00000E86: begin
				q			<=			16'h00D1;
		end
		32'h00000E88: begin
				q			<=			16'h1537;
		end
		32'h00000E8A: begin
				q			<=			16'h0001;
		end
		32'h00000E8C: begin
				q			<=			16'h0693;
		end
		32'h00000E8E: begin
				q			<=			16'hD1C5;
		end
		32'h00000E90: begin
				q			<=			16'h0637;
		end
		32'h00000E92: begin
				q			<=			16'h0001;
		end
		32'h00000E94: begin
				q			<=			16'h0613;
		end
		32'h00000E96: begin
				q			<=			16'hCB86;
		end
		32'h00000E98: begin
				q			<=			16'h0593;
		end
		32'h00000E9A: begin
				q			<=			16'h1000;
		end
		32'h00000E9C: begin
				q			<=			16'h0513;
		end
		32'h00000E9E: begin
				q			<=			16'hD1C5;
		end
		32'h00000EA0: begin
				q			<=			16'h2097;
		end
		32'h00000EA2: begin
				q			<=			16'h0000;
		end
		32'h00000EA4: begin
				q			<=			16'h80E7;
		end
		32'h00000EA6: begin
				q			<=			16'hECC0;
		end
		32'h00000EA8: begin
				q			<=			16'h1793;
		end
		32'h00000EAA: begin
				q			<=			16'h0104;
		end
		32'h00000EAC: begin
				q			<=			16'hCE63;
		end
		32'h00000EAE: begin
				q			<=			16'h2607;
		end
		32'h00000EB0: begin
				q			<=			16'h1737;
		end
		32'h00000EB2: begin
				q			<=			16'h0001;
		end
		32'h00000EB4: begin
				q			<=			16'h0713;
		end
		32'h00000EB6: begin
				q			<=			16'h8E87;
		end
		32'h00000EB8: begin
				q			<=			16'h1793;
		end
		32'h00000EBA: begin
				q			<=			16'h0114;
		end
		32'h00000EBC: begin
				q			<=			16'hCC63;
		end
		32'h00000EBE: begin
				q			<=			16'h2607;
		end
		32'h00000EC0: begin
				q			<=			16'h17B7;
		end
		32'h00000EC2: begin
				q			<=			16'h0001;
		end
		32'h00000EC4: begin
				q			<=			16'h8793;
		end
		32'h00000EC6: begin
				q			<=			16'h8E87;
		end
		32'h00000EC8: begin
				q			<=			16'h1693;
		end
		32'h00000ECA: begin
				q			<=			16'h0124;
		end
		32'h00000ECC: begin
				q			<=			16'hCA63;
		end
		32'h00000ECE: begin
				q			<=			16'h2606;
		end
		32'h00000ED0: begin
				q			<=			16'h1837;
		end
		32'h00000ED2: begin
				q			<=			16'h0001;
		end
		32'h00000ED4: begin
				q			<=			16'h0813;
		end
		32'h00000ED6: begin
				q			<=			16'h8E88;
		end
		32'h00000ED8: begin
				q			<=			16'h1693;
		end
		32'h00000EDA: begin
				q			<=			16'h0134;
		end
		32'h00000EDC: begin
				q			<=			16'hC863;
		end
		32'h00000EDE: begin
				q			<=			16'h2606;
		end
		32'h00000EE0: begin
				q			<=			16'h18B7;
		end
		32'h00000EE2: begin
				q			<=			16'h0001;
		end
		32'h00000EE4: begin
				q			<=			16'h8893;
		end
		32'h00000EE6: begin
				q			<=			16'h8E88;
		end
		32'h00000EE8: begin
				q			<=			16'h1693;
		end
		32'h00000EEA: begin
				q			<=			16'h0144;
		end
		32'h00000EEC: begin
				q			<=			16'hC663;
		end
		32'h00000EEE: begin
				q			<=			16'h2606;
		end
		32'h00000EF0: begin
				q			<=			16'h16B7;
		end
		32'h00000EF2: begin
				q			<=			16'h0001;
		end
		32'h00000EF4: begin
				q			<=			16'h8693;
		end
		32'h00000EF6: begin
				q			<=			16'h8E86;
		end
		32'h00000EF8: begin
				q			<=			16'h5613;
		end
		32'h00000EFA: begin
				q			<=			16'h00A4;
		end
		32'h00000EFC: begin
				q			<=			16'h7613;
		end
		32'h00000EFE: begin
				q			<=			16'h0016;
		end
		32'h00000F00: begin
				q			<=			16'h1263;
		end
		32'h00000F02: begin
				q			<=			16'h2606;
		end
		32'h00000F04: begin
				q			<=			16'h1637;
		end
		32'h00000F06: begin
				q			<=			16'h0001;
		end
		32'h00000F08: begin
				q			<=			16'h0613;
		end
		32'h00000F0A: begin
				q			<=			16'h8E86;
		end
		32'h00000F0C: begin
				q			<=			16'h5593;
		end
		32'h00000F0E: begin
				q			<=			16'h0094;
		end
		32'h00000F10: begin
				q			<=			16'hF593;
		end
		32'h00000F12: begin
				q			<=			16'h0015;
		end
		32'h00000F14: begin
				q			<=			16'h9E63;
		end
		32'h00000F16: begin
				q			<=			16'h2405;
		end
		32'h00000F18: begin
				q			<=			16'h15B7;
		end
		32'h00000F1A: begin
				q			<=			16'h0001;
		end
		32'h00000F1C: begin
				q			<=			16'h8593;
		end
		32'h00000F1E: begin
				q			<=			16'h8E85;
		end
		32'h00000F20: begin
				q			<=			16'h5513;
		end
		32'h00000F22: begin
				q			<=			16'h0084;
		end
		32'h00000F24: begin
				q			<=			16'h7513;
		end
		32'h00000F26: begin
				q			<=			16'h0015;
		end
		32'h00000F28: begin
				q			<=			16'h1A63;
		end
		32'h00000F2A: begin
				q			<=			16'h2405;
		end
		32'h00000F2C: begin
				q			<=			16'h1537;
		end
		32'h00000F2E: begin
				q			<=			16'h0001;
		end
		32'h00000F30: begin
				q			<=			16'h0513;
		end
		32'h00000F32: begin
				q			<=			16'h8E85;
		end
		32'h00000F34: begin
				q			<=			16'h2623;
		end
		32'h00000F36: begin
				q			<=			16'h00A1;
		end
		32'h00000F38: begin
				q			<=			16'h2423;
		end
		32'h00000F3A: begin
				q			<=			16'h00B1;
		end
		32'h00000F3C: begin
				q			<=			16'h2223;
		end
		32'h00000F3E: begin
				q			<=			16'h00C1;
		end
		32'h00000F40: begin
				q			<=			16'h2023;
		end
		32'h00000F42: begin
				q			<=			16'h00D1;
		end
		32'h00000F44: begin
				q			<=			16'h1537;
		end
		32'h00000F46: begin
				q			<=			16'h0001;
		end
		32'h00000F48: begin
				q			<=			16'h0693;
		end
		32'h00000F4A: begin
				q			<=			16'hD1C5;
		end
		32'h00000F4C: begin
				q			<=			16'h0637;
		end
		32'h00000F4E: begin
				q			<=			16'h0001;
		end
		32'h00000F50: begin
				q			<=			16'h0613;
		end
		32'h00000F52: begin
				q			<=			16'hCB86;
		end
		32'h00000F54: begin
				q			<=			16'h0593;
		end
		32'h00000F56: begin
				q			<=			16'h1000;
		end
		32'h00000F58: begin
				q			<=			16'h0513;
		end
		32'h00000F5A: begin
				q			<=			16'hD1C5;
		end
		32'h00000F5C: begin
				q			<=			16'h2097;
		end
		32'h00000F5E: begin
				q			<=			16'h0000;
		end
		32'h00000F60: begin
				q			<=			16'h80E7;
		end
		32'h00000F62: begin
				q			<=			16'hE100;
		end
		32'h00000F64: begin
				q			<=			16'h5793;
		end
		32'h00000F66: begin
				q			<=			16'h0074;
		end
		32'h00000F68: begin
				q			<=			16'hF793;
		end
		32'h00000F6A: begin
				q			<=			16'h0017;
		end
		32'h00000F6C: begin
				q			<=			16'h9E63;
		end
		32'h00000F6E: begin
				q			<=			16'h2007;
		end
		32'h00000F70: begin
				q			<=			16'h1737;
		end
		32'h00000F72: begin
				q			<=			16'h0001;
		end
		32'h00000F74: begin
				q			<=			16'h0713;
		end
		32'h00000F76: begin
				q			<=			16'h8E87;
		end
		32'h00000F78: begin
				q			<=			16'h5793;
		end
		32'h00000F7A: begin
				q			<=			16'h0064;
		end
		32'h00000F7C: begin
				q			<=			16'hF793;
		end
		32'h00000F7E: begin
				q			<=			16'h0017;
		end
		32'h00000F80: begin
				q			<=			16'h9A63;
		end
		32'h00000F82: begin
				q			<=			16'h2007;
		end
		32'h00000F84: begin
				q			<=			16'h17B7;
		end
		32'h00000F86: begin
				q			<=			16'h0001;
		end
		32'h00000F88: begin
				q			<=			16'h8793;
		end
		32'h00000F8A: begin
				q			<=			16'h8E87;
		end
		32'h00000F8C: begin
				q			<=			16'h5693;
		end
		32'h00000F8E: begin
				q			<=			16'h0054;
		end
		32'h00000F90: begin
				q			<=			16'hF693;
		end
		32'h00000F92: begin
				q			<=			16'h0016;
		end
		32'h00000F94: begin
				q			<=			16'h9663;
		end
		32'h00000F96: begin
				q			<=			16'h2006;
		end
		32'h00000F98: begin
				q			<=			16'h1837;
		end
		32'h00000F9A: begin
				q			<=			16'h0001;
		end
		32'h00000F9C: begin
				q			<=			16'h0813;
		end
		32'h00000F9E: begin
				q			<=			16'h8E88;
		end
		32'h00000FA0: begin
				q			<=			16'h5693;
		end
		32'h00000FA2: begin
				q			<=			16'h0044;
		end
		32'h00000FA4: begin
				q			<=			16'hF693;
		end
		32'h00000FA6: begin
				q			<=			16'h0016;
		end
		32'h00000FA8: begin
				q			<=			16'h9263;
		end
		32'h00000FAA: begin
				q			<=			16'h2006;
		end
		32'h00000FAC: begin
				q			<=			16'h18B7;
		end
		32'h00000FAE: begin
				q			<=			16'h0001;
		end
		32'h00000FB0: begin
				q			<=			16'h8893;
		end
		32'h00000FB2: begin
				q			<=			16'h8E88;
		end
		32'h00000FB4: begin
				q			<=			16'h5693;
		end
		32'h00000FB6: begin
				q			<=			16'h0034;
		end
		32'h00000FB8: begin
				q			<=			16'hF693;
		end
		32'h00000FBA: begin
				q			<=			16'h0016;
		end
		32'h00000FBC: begin
				q			<=			16'h9E63;
		end
		32'h00000FBE: begin
				q			<=			16'h1E06;
		end
		32'h00000FC0: begin
				q			<=			16'h16B7;
		end
		32'h00000FC2: begin
				q			<=			16'h0001;
		end
		32'h00000FC4: begin
				q			<=			16'h8693;
		end
		32'h00000FC6: begin
				q			<=			16'h8E86;
		end
		32'h00000FC8: begin
				q			<=			16'h5613;
		end
		32'h00000FCA: begin
				q			<=			16'h0024;
		end
		32'h00000FCC: begin
				q			<=			16'h7613;
		end
		32'h00000FCE: begin
				q			<=			16'h0016;
		end
		32'h00000FD0: begin
				q			<=			16'h1A63;
		end
		32'h00000FD2: begin
				q			<=			16'h1E06;
		end
		32'h00000FD4: begin
				q			<=			16'h1637;
		end
		32'h00000FD6: begin
				q			<=			16'h0001;
		end
		32'h00000FD8: begin
				q			<=			16'h0613;
		end
		32'h00000FDA: begin
				q			<=			16'h8E86;
		end
		32'h00000FDC: begin
				q			<=			16'h5593;
		end
		32'h00000FDE: begin
				q			<=			16'h0014;
		end
		32'h00000FE0: begin
				q			<=			16'hF593;
		end
		32'h00000FE2: begin
				q			<=			16'h0015;
		end
		32'h00000FE4: begin
				q			<=			16'h9663;
		end
		32'h00000FE6: begin
				q			<=			16'h1E05;
		end
		32'h00000FE8: begin
				q			<=			16'h15B7;
		end
		32'h00000FEA: begin
				q			<=			16'h0001;
		end
		32'h00000FEC: begin
				q			<=			16'h8593;
		end
		32'h00000FEE: begin
				q			<=			16'h8E85;
		end
		32'h00000FF0: begin
				q			<=			16'h7413;
		end
		32'h00000FF2: begin
				q			<=			16'h0014;
		end
		32'h00000FF4: begin
				q			<=			16'h1463;
		end
		32'h00000FF6: begin
				q			<=			16'h1E04;
		end
		32'h00000FF8: begin
				q			<=			16'h1537;
		end
		32'h00000FFA: begin
				q			<=			16'h0001;
		end
		32'h00000FFC: begin
				q			<=			16'h0513;
		end
		32'h00000FFE: begin
				q			<=			16'h8E85;
		end
		32'h00001000: begin
				q			<=			16'h2623;
		end
		32'h00001002: begin
				q			<=			16'h00A1;
		end
		32'h00001004: begin
				q			<=			16'h2423;
		end
		32'h00001006: begin
				q			<=			16'h00B1;
		end
		32'h00001008: begin
				q			<=			16'h2223;
		end
		32'h0000100A: begin
				q			<=			16'h00C1;
		end
		32'h0000100C: begin
				q			<=			16'h2023;
		end
		32'h0000100E: begin
				q			<=			16'h00D1;
		end
		32'h00001010: begin
				q			<=			16'h1437;
		end
		32'h00001012: begin
				q			<=			16'h0001;
		end
		32'h00001014: begin
				q			<=			16'h0693;
		end
		32'h00001016: begin
				q			<=			16'hD1C4;
		end
		32'h00001018: begin
				q			<=			16'h0637;
		end
		32'h0000101A: begin
				q			<=			16'h0001;
		end
		32'h0000101C: begin
				q			<=			16'h0613;
		end
		32'h0000101E: begin
				q			<=			16'hCB86;
		end
		32'h00001020: begin
				q			<=			16'h0593;
		end
		32'h00001022: begin
				q			<=			16'h1000;
		end
		32'h00001024: begin
				q			<=			16'h0513;
		end
		32'h00001026: begin
				q			<=			16'hD1C4;
		end
		32'h00001028: begin
				q			<=			16'h2097;
		end
		32'h0000102A: begin
				q			<=			16'h0000;
		end
		32'h0000102C: begin
				q			<=			16'h80E7;
		end
		32'h0000102E: begin
				q			<=			16'hD440;
		end
		32'h00001030: begin
				q			<=			16'h0593;
		end
		32'h00001032: begin
				q			<=			16'h0000;
		end
		32'h00001034: begin
				q			<=			16'h0513;
		end
		32'h00001036: begin
				q			<=			16'hD1C4;
		end
		32'h00001038: begin
				q			<=			16'hF0EF;
		end
		32'h0000103A: begin
				q			<=			16'hB61F;
		end
		32'h0000103C: begin
				q			<=			16'h0513;
		end
		32'h0000103E: begin
				q			<=			16'hD1C4;
		end
		32'h00001040: begin
				q			<=			16'h10EF;
		end
		32'h00001042: begin
				q			<=			16'h5ED0;
		end
		32'h00001044: begin
				q			<=			16'h17B7;
		end
		32'h00001046: begin
				q			<=			16'h0001;
		end
		32'h00001048: begin
				q			<=			16'h8793;
		end
		32'h0000104A: begin
				q			<=			16'hF907;
		end
		32'h0000104C: begin
				q			<=			16'hA703;
		end
		32'h0000104E: begin
				q			<=			16'h0007;
		end
		32'h00001050: begin
				q			<=			16'h0533;
		end
		32'h00001052: begin
				q			<=			16'h00A7;
		end
		32'h00001054: begin
				q			<=			16'hA023;
		end
		32'h00001056: begin
				q			<=			16'h00A7;
		end
		32'h00001058: begin
				q			<=			16'h2083;
		end
		32'h0000105A: begin
				q			<=			16'h01C1;
		end
		32'h0000105C: begin
				q			<=			16'h2403;
		end
		32'h0000105E: begin
				q			<=			16'h0181;
		end
		32'h00001060: begin
				q			<=			16'h0113;
		end
		32'h00001062: begin
				q			<=			16'h0201;
		end
		32'h00001064: begin
				q			<=			16'h8067;
		end
		32'h00001066: begin
				q			<=			16'h0000;
		end
		32'h00001068: begin
				q			<=			16'h16B7;
		end
		32'h0000106A: begin
				q			<=			16'h0001;
		end
		32'h0000106C: begin
				q			<=			16'h8693;
		end
		32'h0000106E: begin
				q			<=			16'h8E46;
		end
		32'h00001070: begin
				q			<=			16'hF06F;
		end
		32'h00001072: begin
				q			<=			16'hCF1F;
		end
		32'h00001074: begin
				q			<=			16'h1737;
		end
		32'h00001076: begin
				q			<=			16'h0001;
		end
		32'h00001078: begin
				q			<=			16'h0713;
		end
		32'h0000107A: begin
				q			<=			16'h8E47;
		end
		32'h0000107C: begin
				q			<=			16'hF06F;
		end
		32'h0000107E: begin
				q			<=			16'hCF5F;
		end
		32'h00001080: begin
				q			<=			16'h17B7;
		end
		32'h00001082: begin
				q			<=			16'h0001;
		end
		32'h00001084: begin
				q			<=			16'h8793;
		end
		32'h00001086: begin
				q			<=			16'h8E47;
		end
		32'h00001088: begin
				q			<=			16'hF06F;
		end
		32'h0000108A: begin
				q			<=			16'hCF9F;
		end
		32'h0000108C: begin
				q			<=			16'h1837;
		end
		32'h0000108E: begin
				q			<=			16'h0001;
		end
		32'h00001090: begin
				q			<=			16'h0813;
		end
		32'h00001092: begin
				q			<=			16'h8E48;
		end
		32'h00001094: begin
				q			<=			16'hF06F;
		end
		32'h00001096: begin
				q			<=			16'hCFDF;
		end
		32'h00001098: begin
				q			<=			16'h18B7;
		end
		32'h0000109A: begin
				q			<=			16'h0001;
		end
		32'h0000109C: begin
				q			<=			16'h8893;
		end
		32'h0000109E: begin
				q			<=			16'h8E48;
		end
		32'h000010A0: begin
				q			<=			16'hF06F;
		end
		32'h000010A2: begin
				q			<=			16'hD01F;
		end
		32'h000010A4: begin
				q			<=			16'h1637;
		end
		32'h000010A6: begin
				q			<=			16'h0001;
		end
		32'h000010A8: begin
				q			<=			16'h0613;
		end
		32'h000010AA: begin
				q			<=			16'h8E46;
		end
		32'h000010AC: begin
				q			<=			16'hF06F;
		end
		32'h000010AE: begin
				q			<=			16'hD05F;
		end
		32'h000010B0: begin
				q			<=			16'h15B7;
		end
		32'h000010B2: begin
				q			<=			16'h0001;
		end
		32'h000010B4: begin
				q			<=			16'h8593;
		end
		32'h000010B6: begin
				q			<=			16'h8E45;
		end
		32'h000010B8: begin
				q			<=			16'hF06F;
		end
		32'h000010BA: begin
				q			<=			16'hD09F;
		end
		32'h000010BC: begin
				q			<=			16'h1537;
		end
		32'h000010BE: begin
				q			<=			16'h0001;
		end
		32'h000010C0: begin
				q			<=			16'h0513;
		end
		32'h000010C2: begin
				q			<=			16'h8E45;
		end
		32'h000010C4: begin
				q			<=			16'hF06F;
		end
		32'h000010C6: begin
				q			<=			16'hD0DF;
		end
		32'h000010C8: begin
				q			<=			16'h1737;
		end
		32'h000010CA: begin
				q			<=			16'h0001;
		end
		32'h000010CC: begin
				q			<=			16'h0713;
		end
		32'h000010CE: begin
				q			<=			16'h8E47;
		end
		32'h000010D0: begin
				q			<=			16'hF06F;
		end
		32'h000010D2: begin
				q			<=			16'hD39F;
		end
		32'h000010D4: begin
				q			<=			16'h17B7;
		end
		32'h000010D6: begin
				q			<=			16'h0001;
		end
		32'h000010D8: begin
				q			<=			16'h8793;
		end
		32'h000010DA: begin
				q			<=			16'h8E47;
		end
		32'h000010DC: begin
				q			<=			16'hF06F;
		end
		32'h000010DE: begin
				q			<=			16'hD3DF;
		end
		32'h000010E0: begin
				q			<=			16'h1837;
		end
		32'h000010E2: begin
				q			<=			16'h0001;
		end
		32'h000010E4: begin
				q			<=			16'h0813;
		end
		32'h000010E6: begin
				q			<=			16'h8E48;
		end
		32'h000010E8: begin
				q			<=			16'hF06F;
		end
		32'h000010EA: begin
				q			<=			16'hD41F;
		end
		32'h000010EC: begin
				q			<=			16'h18B7;
		end
		32'h000010EE: begin
				q			<=			16'h0001;
		end
		32'h000010F0: begin
				q			<=			16'h8893;
		end
		32'h000010F2: begin
				q			<=			16'h8E48;
		end
		32'h000010F4: begin
				q			<=			16'hF06F;
		end
		32'h000010F6: begin
				q			<=			16'hD45F;
		end
		32'h000010F8: begin
				q			<=			16'h16B7;
		end
		32'h000010FA: begin
				q			<=			16'h0001;
		end
		32'h000010FC: begin
				q			<=			16'h8693;
		end
		32'h000010FE: begin
				q			<=			16'h8E46;
		end
		32'h00001100: begin
				q			<=			16'hF06F;
		end
		32'h00001102: begin
				q			<=			16'hD49F;
		end
		32'h00001104: begin
				q			<=			16'h1637;
		end
		32'h00001106: begin
				q			<=			16'h0001;
		end
		32'h00001108: begin
				q			<=			16'h0613;
		end
		32'h0000110A: begin
				q			<=			16'h8E46;
		end
		32'h0000110C: begin
				q			<=			16'hF06F;
		end
		32'h0000110E: begin
				q			<=			16'hD4DF;
		end
		32'h00001110: begin
				q			<=			16'h15B7;
		end
		32'h00001112: begin
				q			<=			16'h0001;
		end
		32'h00001114: begin
				q			<=			16'h8593;
		end
		32'h00001116: begin
				q			<=			16'h8E45;
		end
		32'h00001118: begin
				q			<=			16'hF06F;
		end
		32'h0000111A: begin
				q			<=			16'hD51F;
		end
		32'h0000111C: begin
				q			<=			16'h1537;
		end
		32'h0000111E: begin
				q			<=			16'h0001;
		end
		32'h00001120: begin
				q			<=			16'h0513;
		end
		32'h00001122: begin
				q			<=			16'h8E45;
		end
		32'h00001124: begin
				q			<=			16'hF06F;
		end
		32'h00001126: begin
				q			<=			16'hD55F;
		end
		32'h00001128: begin
				q			<=			16'h1737;
		end
		32'h0000112A: begin
				q			<=			16'h0001;
		end
		32'h0000112C: begin
				q			<=			16'h0713;
		end
		32'h0000112E: begin
				q			<=			16'h8E47;
		end
		32'h00001130: begin
				q			<=			16'hF06F;
		end
		32'h00001132: begin
				q			<=			16'hD89F;
		end
		32'h00001134: begin
				q			<=			16'h17B7;
		end
		32'h00001136: begin
				q			<=			16'h0001;
		end
		32'h00001138: begin
				q			<=			16'h8793;
		end
		32'h0000113A: begin
				q			<=			16'h8E47;
		end
		32'h0000113C: begin
				q			<=			16'hF06F;
		end
		32'h0000113E: begin
				q			<=			16'hD8DF;
		end
		32'h00001140: begin
				q			<=			16'h1837;
		end
		32'h00001142: begin
				q			<=			16'h0001;
		end
		32'h00001144: begin
				q			<=			16'h0813;
		end
		32'h00001146: begin
				q			<=			16'h8E48;
		end
		32'h00001148: begin
				q			<=			16'hF06F;
		end
		32'h0000114A: begin
				q			<=			16'hD91F;
		end
		32'h0000114C: begin
				q			<=			16'h18B7;
		end
		32'h0000114E: begin
				q			<=			16'h0001;
		end
		32'h00001150: begin
				q			<=			16'h8893;
		end
		32'h00001152: begin
				q			<=			16'h8E48;
		end
		32'h00001154: begin
				q			<=			16'hF06F;
		end
		32'h00001156: begin
				q			<=			16'hD95F;
		end
		32'h00001158: begin
				q			<=			16'h16B7;
		end
		32'h0000115A: begin
				q			<=			16'h0001;
		end
		32'h0000115C: begin
				q			<=			16'h8693;
		end
		32'h0000115E: begin
				q			<=			16'h8E46;
		end
		32'h00001160: begin
				q			<=			16'hF06F;
		end
		32'h00001162: begin
				q			<=			16'hD99F;
		end
		32'h00001164: begin
				q			<=			16'h1637;
		end
		32'h00001166: begin
				q			<=			16'h0001;
		end
		32'h00001168: begin
				q			<=			16'h0613;
		end
		32'h0000116A: begin
				q			<=			16'h8E46;
		end
		32'h0000116C: begin
				q			<=			16'hF06F;
		end
		32'h0000116E: begin
				q			<=			16'hDA1F;
		end
		32'h00001170: begin
				q			<=			16'h15B7;
		end
		32'h00001172: begin
				q			<=			16'h0001;
		end
		32'h00001174: begin
				q			<=			16'h8593;
		end
		32'h00001176: begin
				q			<=			16'h8E45;
		end
		32'h00001178: begin
				q			<=			16'hF06F;
		end
		32'h0000117A: begin
				q			<=			16'hDA9F;
		end
		32'h0000117C: begin
				q			<=			16'h1537;
		end
		32'h0000117E: begin
				q			<=			16'h0001;
		end
		32'h00001180: begin
				q			<=			16'h0513;
		end
		32'h00001182: begin
				q			<=			16'h8E45;
		end
		32'h00001184: begin
				q			<=			16'hF06F;
		end
		32'h00001186: begin
				q			<=			16'hDB1F;
		end
		32'h00001188: begin
				q			<=			16'h1737;
		end
		32'h0000118A: begin
				q			<=			16'h0001;
		end
		32'h0000118C: begin
				q			<=			16'h0713;
		end
		32'h0000118E: begin
				q			<=			16'h8E47;
		end
		32'h00001190: begin
				q			<=			16'hF06F;
		end
		32'h00001192: begin
				q			<=			16'hDE9F;
		end
		32'h00001194: begin
				q			<=			16'h17B7;
		end
		32'h00001196: begin
				q			<=			16'h0001;
		end
		32'h00001198: begin
				q			<=			16'h8793;
		end
		32'h0000119A: begin
				q			<=			16'h8E47;
		end
		32'h0000119C: begin
				q			<=			16'hF06F;
		end
		32'h0000119E: begin
				q			<=			16'hDF1F;
		end
		32'h000011A0: begin
				q			<=			16'h1837;
		end
		32'h000011A2: begin
				q			<=			16'h0001;
		end
		32'h000011A4: begin
				q			<=			16'h0813;
		end
		32'h000011A6: begin
				q			<=			16'h8E48;
		end
		32'h000011A8: begin
				q			<=			16'hF06F;
		end
		32'h000011AA: begin
				q			<=			16'hDF9F;
		end
		32'h000011AC: begin
				q			<=			16'h18B7;
		end
		32'h000011AE: begin
				q			<=			16'h0001;
		end
		32'h000011B0: begin
				q			<=			16'h8893;
		end
		32'h000011B2: begin
				q			<=			16'h8E48;
		end
		32'h000011B4: begin
				q			<=			16'hF06F;
		end
		32'h000011B6: begin
				q			<=			16'hE01F;
		end
		32'h000011B8: begin
				q			<=			16'h16B7;
		end
		32'h000011BA: begin
				q			<=			16'h0001;
		end
		32'h000011BC: begin
				q			<=			16'h8693;
		end
		32'h000011BE: begin
				q			<=			16'h8E46;
		end
		32'h000011C0: begin
				q			<=			16'hF06F;
		end
		32'h000011C2: begin
				q			<=			16'hE09F;
		end
		32'h000011C4: begin
				q			<=			16'h1637;
		end
		32'h000011C6: begin
				q			<=			16'h0001;
		end
		32'h000011C8: begin
				q			<=			16'h0613;
		end
		32'h000011CA: begin
				q			<=			16'h8E46;
		end
		32'h000011CC: begin
				q			<=			16'hF06F;
		end
		32'h000011CE: begin
				q			<=			16'hE11F;
		end
		32'h000011D0: begin
				q			<=			16'h15B7;
		end
		32'h000011D2: begin
				q			<=			16'h0001;
		end
		32'h000011D4: begin
				q			<=			16'h8593;
		end
		32'h000011D6: begin
				q			<=			16'h8E45;
		end
		32'h000011D8: begin
				q			<=			16'hF06F;
		end
		32'h000011DA: begin
				q			<=			16'hE19F;
		end
		32'h000011DC: begin
				q			<=			16'h1537;
		end
		32'h000011DE: begin
				q			<=			16'h0001;
		end
		32'h000011E0: begin
				q			<=			16'h0513;
		end
		32'h000011E2: begin
				q			<=			16'h8E45;
		end
		32'h000011E4: begin
				q			<=			16'hF06F;
		end
		32'h000011E6: begin
				q			<=			16'hE1DF;
		end
		32'h000011E8: begin
				q			<=			16'h0000;
		end
		32'h000011EA: begin
				q			<=			16'h0000;
		end
		32'h000011EC: begin
				q			<=			16'h0113;
		end
		32'h000011EE: begin
				q			<=			16'hFF01;
		end
		32'h000011F0: begin
				q			<=			16'h2623;
		end
		32'h000011F2: begin
				q			<=			16'h0011;
		end
		32'h000011F4: begin
				q			<=			16'h2423;
		end
		32'h000011F6: begin
				q			<=			16'h0081;
		end
		32'h000011F8: begin
				q			<=			16'h1693;
		end
		32'h000011FA: begin
				q			<=			16'h0105;
		end
		32'h000011FC: begin
				q			<=			16'hD693;
		end
		32'h000011FE: begin
				q			<=			16'h0106;
		end
		32'h00001200: begin
				q			<=			16'h0637;
		end
		32'h00001202: begin
				q			<=			16'h0001;
		end
		32'h00001204: begin
				q			<=			16'h0613;
		end
		32'h00001206: begin
				q			<=			16'hCCC6;
		end
		32'h00001208: begin
				q			<=			16'h0593;
		end
		32'h0000120A: begin
				q			<=			16'h1000;
		end
		32'h0000120C: begin
				q			<=			16'h1437;
		end
		32'h0000120E: begin
				q			<=			16'h0001;
		end
		32'h00001210: begin
				q			<=			16'h0513;
		end
		32'h00001212: begin
				q			<=			16'hD1C4;
		end
		32'h00001214: begin
				q			<=			16'h2097;
		end
		32'h00001216: begin
				q			<=			16'h0000;
		end
		32'h00001218: begin
				q			<=			16'h80E7;
		end
		32'h0000121A: begin
				q			<=			16'hB580;
		end
		32'h0000121C: begin
				q			<=			16'h0593;
		end
		32'h0000121E: begin
				q			<=			16'h0000;
		end
		32'h00001220: begin
				q			<=			16'h0513;
		end
		32'h00001222: begin
				q			<=			16'hD1C4;
		end
		32'h00001224: begin
				q			<=			16'hF0EF;
		end
		32'h00001226: begin
				q			<=			16'h975F;
		end
		32'h00001228: begin
				q			<=			16'h0513;
		end
		32'h0000122A: begin
				q			<=			16'hD1C4;
		end
		32'h0000122C: begin
				q			<=			16'h10EF;
		end
		32'h0000122E: begin
				q			<=			16'h4010;
		end
		32'h00001230: begin
				q			<=			16'h17B7;
		end
		32'h00001232: begin
				q			<=			16'h0001;
		end
		32'h00001234: begin
				q			<=			16'h8793;
		end
		32'h00001236: begin
				q			<=			16'hF907;
		end
		32'h00001238: begin
				q			<=			16'hA703;
		end
		32'h0000123A: begin
				q			<=			16'h0007;
		end
		32'h0000123C: begin
				q			<=			16'h0533;
		end
		32'h0000123E: begin
				q			<=			16'h00A7;
		end
		32'h00001240: begin
				q			<=			16'hA023;
		end
		32'h00001242: begin
				q			<=			16'h00A7;
		end
		32'h00001244: begin
				q			<=			16'h2083;
		end
		32'h00001246: begin
				q			<=			16'h00C1;
		end
		32'h00001248: begin
				q			<=			16'h2403;
		end
		32'h0000124A: begin
				q			<=			16'h0081;
		end
		32'h0000124C: begin
				q			<=			16'h0113;
		end
		32'h0000124E: begin
				q			<=			16'h0101;
		end
		32'h00001250: begin
				q			<=			16'h8067;
		end
		32'h00001252: begin
				q			<=			16'h0000;
		end
		32'h00001254: begin
				q			<=			16'h0000;
		end
		32'h00001256: begin
				q			<=			16'h0000;
		end
		32'h00001258: begin
				q			<=			16'h4783;
		end
		32'h0000125A: begin
				q			<=			16'h0005;
		end
		32'h0000125C: begin
				q			<=			16'hF793;
		end
		32'h0000125E: begin
				q			<=			16'h0DF7;
		end
		32'h00001260: begin
				q			<=			16'h8263;
		end
		32'h00001262: begin
				q			<=			16'h0207;
		end
		32'h00001264: begin
				q			<=			16'h0713;
		end
		32'h00001266: begin
				q			<=			16'h0015;
		end
		32'h00001268: begin
				q			<=			16'h0513;
		end
		32'h0000126A: begin
				q			<=			16'h0000;
		end
		32'h0000126C: begin
				q			<=			16'h0513;
		end
		32'h0000126E: begin
				q			<=			16'h0015;
		end
		32'h00001270: begin
				q			<=			16'h4783;
		end
		32'h00001272: begin
				q			<=			16'h0007;
		end
		32'h00001274: begin
				q			<=			16'hF793;
		end
		32'h00001276: begin
				q			<=			16'h0DF7;
		end
		32'h00001278: begin
				q			<=			16'h0713;
		end
		32'h0000127A: begin
				q			<=			16'h0017;
		end
		32'h0000127C: begin
				q			<=			16'h98E3;
		end
		32'h0000127E: begin
				q			<=			16'hFE07;
		end
		32'h00001280: begin
				q			<=			16'h8067;
		end
		32'h00001282: begin
				q			<=			16'h0000;
		end
		32'h00001284: begin
				q			<=			16'h0513;
		end
		32'h00001286: begin
				q			<=			16'h0000;
		end
		32'h00001288: begin
				q			<=			16'h8067;
		end
		32'h0000128A: begin
				q			<=			16'h0000;
		end
		32'h0000128C: begin
				q			<=			16'h0000;
		end
		32'h0000128E: begin
				q			<=			16'h0000;
		end
		32'h00001290: begin
				q			<=			16'h17B7;
		end
		32'h00001292: begin
				q			<=			16'h0001;
		end
		32'h00001294: begin
				q			<=			16'hAA23;
		end
		32'h00001296: begin
				q			<=			16'hF8A7;
		end
		32'h00001298: begin
				q			<=			16'h8067;
		end
		32'h0000129A: begin
				q			<=			16'h0000;
		end
		32'h0000129C: begin
				q			<=			16'h0000;
		end
		32'h0000129E: begin
				q			<=			16'h0000;
		end
		32'h000012A0: begin
				q			<=			16'h17B7;
		end
		32'h000012A2: begin
				q			<=			16'h0001;
		end
		32'h000012A4: begin
				q			<=			16'hA503;
		end
		32'h000012A6: begin
				q			<=			16'hF947;
		end
		32'h000012A8: begin
				q			<=			16'h8067;
		end
		32'h000012AA: begin
				q			<=			16'h0000;
		end
		32'h000012AC: begin
				q			<=			16'h0000;
		end
		32'h000012AE: begin
				q			<=			16'h0000;
		end
		32'h000012B0: begin
				q			<=			16'h0113;
		end
		32'h000012B2: begin
				q			<=			16'hFF01;
		end
		32'h000012B4: begin
				q			<=			16'h2623;
		end
		32'h000012B6: begin
				q			<=			16'h0011;
		end
		32'h000012B8: begin
				q			<=			16'h2423;
		end
		32'h000012BA: begin
				q			<=			16'h0081;
		end
		32'h000012BC: begin
				q			<=			16'h0693;
		end
		32'h000012BE: begin
				q			<=			16'h0005;
		end
		32'h000012C0: begin
				q			<=			16'h0637;
		end
		32'h000012C2: begin
				q			<=			16'h0001;
		end
		32'h000012C4: begin
				q			<=			16'h0613;
		end
		32'h000012C6: begin
				q			<=			16'hCE86;
		end
		32'h000012C8: begin
				q			<=			16'h0593;
		end
		32'h000012CA: begin
				q			<=			16'h1000;
		end
		32'h000012CC: begin
				q			<=			16'h1437;
		end
		32'h000012CE: begin
				q			<=			16'h0001;
		end
		32'h000012D0: begin
				q			<=			16'h0513;
		end
		32'h000012D2: begin
				q			<=			16'hD1C4;
		end
		32'h000012D4: begin
				q			<=			16'h2097;
		end
		32'h000012D6: begin
				q			<=			16'h0000;
		end
		32'h000012D8: begin
				q			<=			16'h80E7;
		end
		32'h000012DA: begin
				q			<=			16'hA980;
		end
		32'h000012DC: begin
				q			<=			16'h0593;
		end
		32'h000012DE: begin
				q			<=			16'h0010;
		end
		32'h000012E0: begin
				q			<=			16'h0513;
		end
		32'h000012E2: begin
				q			<=			16'hD1C4;
		end
		32'h000012E4: begin
				q			<=			16'hF0EF;
		end
		32'h000012E6: begin
				q			<=			16'h8B5F;
		end
		32'h000012E8: begin
				q			<=			16'h006F;
		end
		32'h000012EA: begin
				q			<=			16'h0000;
		end
		32'h000012EC: begin
				q			<=			16'h0000;
		end
		32'h000012EE: begin
				q			<=			16'h0000;
		end
		32'h000012F0: begin
				q			<=			16'h0113;
		end
		32'h000012F2: begin
				q			<=			16'hFF01;
		end
		32'h000012F4: begin
				q			<=			16'h2623;
		end
		32'h000012F6: begin
				q			<=			16'h0011;
		end
		32'h000012F8: begin
				q			<=			16'h17B7;
		end
		32'h000012FA: begin
				q			<=			16'h0001;
		end
		32'h000012FC: begin
				q			<=			16'h8793;
		end
		32'h000012FE: begin
				q			<=			16'hF947;
		end
		32'h00001300: begin
				q			<=			16'hA683;
		end
		32'h00001302: begin
				q			<=			16'h0007;
		end
		32'h00001304: begin
				q			<=			16'h0713;
		end
		32'h00001306: begin
				q			<=			16'h0040;
		end
		32'h00001308: begin
				q			<=			16'h6463;
		end
		32'h0000130A: begin
				q			<=			16'h08D7;
		end
		32'h0000130C: begin
				q			<=			16'h9793;
		end
		32'h0000130E: begin
				q			<=			16'h0026;
		end
		32'h00001310: begin
				q			<=			16'h0737;
		end
		32'h00001312: begin
				q			<=			16'h0001;
		end
		32'h00001314: begin
				q			<=			16'h0713;
		end
		32'h00001316: begin
				q			<=			16'hCD47;
		end
		32'h00001318: begin
				q			<=			16'h87B3;
		end
		32'h0000131A: begin
				q			<=			16'h00E7;
		end
		32'h0000131C: begin
				q			<=			16'hA783;
		end
		32'h0000131E: begin
				q			<=			16'h0007;
		end
		32'h00001320: begin
				q			<=			16'h8067;
		end
		32'h00001322: begin
				q			<=			16'h0007;
		end
		32'h00001324: begin
				q			<=			16'h0593;
		end
		32'h00001326: begin
				q			<=			16'h0010;
		end
		32'h00001328: begin
				q			<=			16'h0537;
		end
		32'h0000132A: begin
				q			<=			16'h0001;
		end
		32'h0000132C: begin
				q			<=			16'h0513;
		end
		32'h0000132E: begin
				q			<=			16'hCF85;
		end
		32'h00001330: begin
				q			<=			16'hF0EF;
		end
		32'h00001332: begin
				q			<=			16'h869F;
		end
		32'h00001334: begin
				q			<=			16'h2083;
		end
		32'h00001336: begin
				q			<=			16'h00C1;
		end
		32'h00001338: begin
				q			<=			16'h0113;
		end
		32'h0000133A: begin
				q			<=			16'h0101;
		end
		32'h0000133C: begin
				q			<=			16'h8067;
		end
		32'h0000133E: begin
				q			<=			16'h0000;
		end
		32'h00001340: begin
				q			<=			16'h0593;
		end
		32'h00001342: begin
				q			<=			16'h0010;
		end
		32'h00001344: begin
				q			<=			16'h0537;
		end
		32'h00001346: begin
				q			<=			16'h0001;
		end
		32'h00001348: begin
				q			<=			16'h0513;
		end
		32'h0000134A: begin
				q			<=			16'hD045;
		end
		32'h0000134C: begin
				q			<=			16'hF0EF;
		end
		32'h0000134E: begin
				q			<=			16'h84DF;
		end
		32'h00001350: begin
				q			<=			16'hF06F;
		end
		32'h00001352: begin
				q			<=			16'hFE5F;
		end
		32'h00001354: begin
				q			<=			16'h0593;
		end
		32'h00001356: begin
				q			<=			16'h0010;
		end
		32'h00001358: begin
				q			<=			16'h0537;
		end
		32'h0000135A: begin
				q			<=			16'h0001;
		end
		32'h0000135C: begin
				q			<=			16'h0513;
		end
		32'h0000135E: begin
				q			<=			16'hD185;
		end
		32'h00001360: begin
				q			<=			16'hF0EF;
		end
		32'h00001362: begin
				q			<=			16'h839F;
		end
		32'h00001364: begin
				q			<=			16'hF06F;
		end
		32'h00001366: begin
				q			<=			16'hFD1F;
		end
		32'h00001368: begin
				q			<=			16'h0593;
		end
		32'h0000136A: begin
				q			<=			16'h0010;
		end
		32'h0000136C: begin
				q			<=			16'h0537;
		end
		32'h0000136E: begin
				q			<=			16'h0001;
		end
		32'h00001370: begin
				q			<=			16'h0513;
		end
		32'h00001372: begin
				q			<=			16'hD285;
		end
		32'h00001374: begin
				q			<=			16'hF0EF;
		end
		32'h00001376: begin
				q			<=			16'h825F;
		end
		32'h00001378: begin
				q			<=			16'hF06F;
		end
		32'h0000137A: begin
				q			<=			16'hFBDF;
		end
		32'h0000137C: begin
				q			<=			16'h0593;
		end
		32'h0000137E: begin
				q			<=			16'h0010;
		end
		32'h00001380: begin
				q			<=			16'h0537;
		end
		32'h00001382: begin
				q			<=			16'h0001;
		end
		32'h00001384: begin
				q			<=			16'h0513;
		end
		32'h00001386: begin
				q			<=			16'hD3C5;
		end
		32'h00001388: begin
				q			<=			16'hF0EF;
		end
		32'h0000138A: begin
				q			<=			16'h811F;
		end
		32'h0000138C: begin
				q			<=			16'hF06F;
		end
		32'h0000138E: begin
				q			<=			16'hFA9F;
		end
		32'h00001390: begin
				q			<=			16'h0593;
		end
		32'h00001392: begin
				q			<=			16'h0010;
		end
		32'h00001394: begin
				q			<=			16'h0537;
		end
		32'h00001396: begin
				q			<=			16'h0001;
		end
		32'h00001398: begin
				q			<=			16'h0513;
		end
		32'h0000139A: begin
				q			<=			16'hD4C5;
		end
		32'h0000139C: begin
				q			<=			16'hF0EF;
		end
		32'h0000139E: begin
				q			<=			16'hFFCF;
		end
		32'h000013A0: begin
				q			<=			16'hF06F;
		end
		32'h000013A2: begin
				q			<=			16'hF95F;
		end
		32'h000013A4: begin
				q			<=			16'h0000;
		end
		32'h000013A6: begin
				q			<=			16'h0000;
		end
		32'h000013A8: begin
				q			<=			16'h0113;
		end
		32'h000013AA: begin
				q			<=			16'hFF01;
		end
		32'h000013AC: begin
				q			<=			16'h2623;
		end
		32'h000013AE: begin
				q			<=			16'h0081;
		end
		32'h000013B0: begin
				q			<=			16'h0413;
		end
		32'h000013B2: begin
				q			<=			16'h0101;
		end
		32'h000013B4: begin
				q			<=			16'h0793;
		end
		32'h000013B6: begin
				q			<=			16'h0030;
		end
		32'h000013B8: begin
				q			<=			16'h0693;
		end
		32'h000013BA: begin
				q			<=			16'h0080;
		end
		32'h000013BC: begin
				q			<=			16'hFA63;
		end
		32'h000013BE: begin
				q			<=			16'h00A7;
		end
		32'h000013C0: begin
				q			<=			16'h06B3;
		end
		32'h000013C2: begin
				q			<=			16'h40A0;
		end
		32'h000013C4: begin
				q			<=			16'hF693;
		end
		32'h000013C6: begin
				q			<=			16'h0036;
		end
		32'h000013C8: begin
				q			<=			16'h0513;
		end
		32'h000013CA: begin
				q			<=			16'h0045;
		end
		32'h000013CC: begin
				q			<=			16'h86B3;
		end
		32'h000013CE: begin
				q			<=			16'h00A6;
		end
		32'h000013D0: begin
				q			<=			16'h17B7;
		end
		32'h000013D2: begin
				q			<=			16'h0001;
		end
		32'h000013D4: begin
				q			<=			16'hA783;
		end
		32'h000013D6: begin
				q			<=			16'hE1C7;
		end
		32'h000013D8: begin
				q			<=			16'h8C63;
		end
		32'h000013DA: begin
				q			<=			16'h0A07;
		end
		32'h000013DC: begin
				q			<=			16'hA703;
		end
		32'h000013DE: begin
				q			<=			16'h0007;
		end
		32'h000013E0: begin
				q			<=			16'h1637;
		end
		32'h000013E2: begin
				q			<=			16'h0001;
		end
		32'h000013E4: begin
				q			<=			16'h0613;
		end
		32'h000013E6: begin
				q			<=			16'hE1C6;
		end
		32'h000013E8: begin
				q			<=			16'h6863;
		end
		32'h000013EA: begin
				q			<=			16'h08D7;
		end
		32'h000013EC: begin
				q			<=			16'h8513;
		end
		32'h000013EE: begin
				q			<=			16'h0007;
		end
		32'h000013F0: begin
				q			<=			16'h1637;
		end
		32'h000013F2: begin
				q			<=			16'h0001;
		end
		32'h000013F4: begin
				q			<=			16'h0613;
		end
		32'h000013F6: begin
				q			<=			16'hE1C6;
		end
		32'h000013F8: begin
				q			<=			16'h8793;
		end
		32'h000013FA: begin
				q			<=			16'h0086;
		end
		32'h000013FC: begin
				q			<=			16'h6263;
		end
		32'h000013FE: begin
				q			<=			16'h02F7;
		end
		32'h00001400: begin
				q			<=			16'h2583;
		end
		32'h00001402: begin
				q			<=			16'h0045;
		end
		32'h00001404: begin
				q			<=			16'h07B3;
		end
		32'h00001406: begin
				q			<=			16'h00D5;
		end
		32'h00001408: begin
				q			<=			16'h2023;
		end
		32'h0000140A: begin
				q			<=			16'h00F6;
		end
		32'h0000140C: begin
				q			<=			16'h0733;
		end
		32'h0000140E: begin
				q			<=			16'h40D7;
		end
		32'h00001410: begin
				q			<=			16'hA023;
		end
		32'h00001412: begin
				q			<=			16'h00E7;
		end
		32'h00001414: begin
				q			<=			16'h2783;
		end
		32'h00001416: begin
				q			<=			16'h0006;
		end
		32'h00001418: begin
				q			<=			16'hA223;
		end
		32'h0000141A: begin
				q			<=			16'h00B7;
		end
		32'h0000141C: begin
				q			<=			16'h006F;
		end
		32'h0000141E: begin
				q			<=			16'h0940;
		end
		32'h00001420: begin
				q			<=			16'h2783;
		end
		32'h00001422: begin
				q			<=			16'h0045;
		end
		32'h00001424: begin
				q			<=			16'h2023;
		end
		32'h00001426: begin
				q			<=			16'h00F6;
		end
		32'h00001428: begin
				q			<=			16'h0513;
		end
		32'h0000142A: begin
				q			<=			16'h0045;
		end
		32'h0000142C: begin
				q			<=			16'h006F;
		end
		32'h0000142E: begin
				q			<=			16'h08C0;
		end
		32'h00001430: begin
				q			<=			16'h05B3;
		end
		32'h00001432: begin
				q			<=			16'h40A4;
		end
		32'h00001434: begin
				q			<=			16'h8593;
		end
		32'h00001436: begin
				q			<=			16'hFE05;
		end
		32'h00001438: begin
				q			<=			16'h8733;
		end
		32'h0000143A: begin
				q			<=			16'h40E6;
		end
		32'h0000143C: begin
				q			<=			16'hEE63;
		end
		32'h0000143E: begin
				q			<=			16'h00E5;
		end
		32'h00001440: begin
				q			<=			16'h2023;
		end
		32'h00001442: begin
				q			<=			16'h0006;
		end
		32'h00001444: begin
				q			<=			16'h8833;
		end
		32'h00001446: begin
				q			<=			16'h00D7;
		end
		32'h00001448: begin
				q			<=			16'h1737;
		end
		32'h0000144A: begin
				q			<=			16'h0001;
		end
		32'h0000144C: begin
				q			<=			16'h2623;
		end
		32'h0000144E: begin
				q			<=			16'h8F07;
		end
		32'h00001450: begin
				q			<=			16'h8513;
		end
		32'h00001452: begin
				q			<=			16'h0007;
		end
		32'h00001454: begin
				q			<=			16'h006F;
		end
		32'h00001456: begin
				q			<=			16'h05C0;
		end
		32'h00001458: begin
				q			<=			16'h0513;
		end
		32'h0000145A: begin
				q			<=			16'h0000;
		end
		32'h0000145C: begin
				q			<=			16'h006F;
		end
		32'h0000145E: begin
				q			<=			16'h05C0;
		end
		32'h00001460: begin
				q			<=			16'h0513;
		end
		32'h00001462: begin
				q			<=			16'h0000;
		end
		32'h00001464: begin
				q			<=			16'h006F;
		end
		32'h00001466: begin
				q			<=			16'h0540;
		end
		32'h00001468: begin
				q			<=			16'h8613;
		end
		32'h0000146A: begin
				q			<=			16'h0047;
		end
		32'h0000146C: begin
				q			<=			16'h2703;
		end
		32'h0000146E: begin
				q			<=			16'h0005;
		end
		32'h00001470: begin
				q			<=			16'h0793;
		end
		32'h00001472: begin
				q			<=			16'h0005;
		end
		32'h00001474: begin
				q			<=			16'h72E3;
		end
		32'h00001476: begin
				q			<=			16'hF8D7;
		end
		32'h00001478: begin
				q			<=			16'hA503;
		end
		32'h0000147A: begin
				q			<=			16'h0047;
		end
		32'h0000147C: begin
				q			<=			16'h16E3;
		end
		32'h0000147E: begin
				q			<=			16'hFE05;
		end
		32'h00001480: begin
				q			<=			16'h85B3;
		end
		32'h00001482: begin
				q			<=			16'h00E7;
		end
		32'h00001484: begin
				q			<=			16'h1537;
		end
		32'h00001486: begin
				q			<=			16'h0001;
		end
		32'h00001488: begin
				q			<=			16'h2503;
		end
		32'h0000148A: begin
				q			<=			16'h8EC5;
		end
		32'h0000148C: begin
				q			<=			16'h02E3;
		end
		32'h0000148E: begin
				q			<=			16'hFAB5;
		end
		32'h00001490: begin
				q			<=			16'h17B7;
		end
		32'h00001492: begin
				q			<=			16'h0001;
		end
		32'h00001494: begin
				q			<=			16'hA503;
		end
		32'h00001496: begin
				q			<=			16'h8EC7;
		end
		32'h00001498: begin
				q			<=			16'h07B3;
		end
		32'h0000149A: begin
				q			<=			16'h40A4;
		end
		32'h0000149C: begin
				q			<=			16'h8793;
		end
		32'h0000149E: begin
				q			<=			16'hFE07;
		end
		32'h000014A0: begin
				q			<=			16'hE0E3;
		end
		32'h000014A2: begin
				q			<=			16'hFCD7;
		end
		32'h000014A4: begin
				q			<=			16'h07B3;
		end
		32'h000014A6: begin
				q			<=			16'h00D5;
		end
		32'h000014A8: begin
				q			<=			16'h1737;
		end
		32'h000014AA: begin
				q			<=			16'h0001;
		end
		32'h000014AC: begin
				q			<=			16'h2623;
		end
		32'h000014AE: begin
				q			<=			16'h8EF7;
		end
		32'h000014B0: begin
				q			<=			16'h2023;
		end
		32'h000014B2: begin
				q			<=			16'h00D5;
		end
		32'h000014B4: begin
				q			<=			16'h0513;
		end
		32'h000014B6: begin
				q			<=			16'h0045;
		end
		32'h000014B8: begin
				q			<=			16'h2403;
		end
		32'h000014BA: begin
				q			<=			16'h00C1;
		end
		32'h000014BC: begin
				q			<=			16'h0113;
		end
		32'h000014BE: begin
				q			<=			16'h0101;
		end
		32'h000014C0: begin
				q			<=			16'h8067;
		end
		32'h000014C2: begin
				q			<=			16'h0000;
		end
		32'h000014C4: begin
				q			<=			16'h0000;
		end
		32'h000014C6: begin
				q			<=			16'h0000;
		end
		32'h000014C8: begin
				q			<=			16'h0C63;
		end
		32'h000014CA: begin
				q			<=			16'h0405;
		end
		32'h000014CC: begin
				q			<=			16'h0713;
		end
		32'h000014CE: begin
				q			<=			16'hFFC5;
		end
		32'h000014D0: begin
				q			<=			16'h17B7;
		end
		32'h000014D2: begin
				q			<=			16'h0001;
		end
		32'h000014D4: begin
				q			<=			16'hA783;
		end
		32'h000014D6: begin
				q			<=			16'hE1C7;
		end
		32'h000014D8: begin
				q			<=			16'h8263;
		end
		32'h000014DA: begin
				q			<=			16'h0A07;
		end
		32'h000014DC: begin
				q			<=			16'hA603;
		end
		32'h000014DE: begin
				q			<=			16'h0007;
		end
		32'h000014E0: begin
				q			<=			16'h05B3;
		end
		32'h000014E2: begin
				q			<=			16'h00F6;
		end
		32'h000014E4: begin
				q			<=			16'h0063;
		end
		32'h000014E6: begin
				q			<=			16'h04B7;
		end
		32'h000014E8: begin
				q			<=			16'h2303;
		end
		32'h000014EA: begin
				q			<=			16'hFFC5;
		end
		32'h000014EC: begin
				q			<=			16'h0833;
		end
		32'h000014EE: begin
				q			<=			16'h0067;
		end
		32'h000014F0: begin
				q			<=			16'h8663;
		end
		32'h000014F2: begin
				q			<=			16'h0707;
		end
		32'h000014F4: begin
				q			<=			16'h6A63;
		end
		32'h000014F6: begin
				q			<=			16'h08F7;
		end
		32'h000014F8: begin
				q			<=			16'h8893;
		end
		32'h000014FA: begin
				q			<=			16'h0047;
		end
		32'h000014FC: begin
				q			<=			16'hA783;
		end
		32'h000014FE: begin
				q			<=			16'h0047;
		end
		32'h00001500: begin
				q			<=			16'h8C63;
		end
		32'h00001502: begin
				q			<=			16'h0007;
		end
		32'h00001504: begin
				q			<=			16'hA603;
		end
		32'h00001506: begin
				q			<=			16'h0007;
		end
		32'h00001508: begin
				q			<=			16'h05B3;
		end
		32'h0000150A: begin
				q			<=			16'h00F6;
		end
		32'h0000150C: begin
				q			<=			16'h0C63;
		end
		32'h0000150E: begin
				q			<=			16'h00B7;
		end
		32'h00001510: begin
				q			<=			16'h8A63;
		end
		32'h00001512: begin
				q			<=			16'h0507;
		end
		32'h00001514: begin
				q			<=			16'h72E3;
		end
		32'h00001516: begin
				q			<=			16'hFEF7;
		end
		32'h00001518: begin
				q			<=			16'h2223;
		end
		32'h0000151A: begin
				q			<=			16'h00F7;
		end
		32'h0000151C: begin
				q			<=			16'hA023;
		end
		32'h0000151E: begin
				q			<=			16'h00E8;
		end
		32'h00001520: begin
				q			<=			16'h8067;
		end
		32'h00001522: begin
				q			<=			16'h0000;
		end
		32'h00001524: begin
				q			<=			16'h2683;
		end
		32'h00001526: begin
				q			<=			16'hFFC5;
		end
		32'h00001528: begin
				q			<=			16'h0633;
		end
		32'h0000152A: begin
				q			<=			16'h00D6;
		end
		32'h0000152C: begin
				q			<=			16'hA023;
		end
		32'h0000152E: begin
				q			<=			16'h00C7;
		end
		32'h00001530: begin
				q			<=			16'hA683;
		end
		32'h00001532: begin
				q			<=			16'h0047;
		end
		32'h00001534: begin
				q			<=			16'h86E3;
		end
		32'h00001536: begin
				q			<=			16'hFE06;
		end
		32'h00001538: begin
				q			<=			16'h2583;
		end
		32'h0000153A: begin
				q			<=			16'hFFC5;
		end
		32'h0000153C: begin
				q			<=			16'h0733;
		end
		32'h0000153E: begin
				q			<=			16'h00B7;
		end
		32'h00001540: begin
				q			<=			16'h90E3;
		end
		32'h00001542: begin
				q			<=			16'hFEE6;
		end
		32'h00001544: begin
				q			<=			16'hA703;
		end
		32'h00001546: begin
				q			<=			16'h0006;
		end
		32'h00001548: begin
				q			<=			16'h0633;
		end
		32'h0000154A: begin
				q			<=			16'h00C7;
		end
		32'h0000154C: begin
				q			<=			16'hA023;
		end
		32'h0000154E: begin
				q			<=			16'h00C7;
		end
		32'h00001550: begin
				q			<=			16'hA703;
		end
		32'h00001552: begin
				q			<=			16'h0046;
		end
		32'h00001554: begin
				q			<=			16'hA223;
		end
		32'h00001556: begin
				q			<=			16'h00E7;
		end
		32'h00001558: begin
				q			<=			16'h8067;
		end
		32'h0000155A: begin
				q			<=			16'h0000;
		end
		32'h0000155C: begin
				q			<=			16'h18B7;
		end
		32'h0000155E: begin
				q			<=			16'h0001;
		end
		32'h00001560: begin
				q			<=			16'h8893;
		end
		32'h00001562: begin
				q			<=			16'hE1C8;
		end
		32'h00001564: begin
				q			<=			16'h0633;
		end
		32'h00001566: begin
				q			<=			16'h00C3;
		end
		32'h00001568: begin
				q			<=			16'h2E23;
		end
		32'h0000156A: begin
				q			<=			16'hFEC5;
		end
		32'h0000156C: begin
				q			<=			16'hA783;
		end
		32'h0000156E: begin
				q			<=			16'h0047;
		end
		32'h00001570: begin
				q			<=			16'h2223;
		end
		32'h00001572: begin
				q			<=			16'h00F7;
		end
		32'h00001574: begin
				q			<=			16'hA023;
		end
		32'h00001576: begin
				q			<=			16'h00E8;
		end
		32'h00001578: begin
				q			<=			16'h8067;
		end
		32'h0000157A: begin
				q			<=			16'h0000;
		end
		32'h0000157C: begin
				q			<=			16'h18B7;
		end
		32'h0000157E: begin
				q			<=			16'h0001;
		end
		32'h00001580: begin
				q			<=			16'h8893;
		end
		32'h00001582: begin
				q			<=			16'hE1C8;
		end
		32'h00001584: begin
				q			<=			16'hF06F;
		end
		32'h00001586: begin
				q			<=			16'hF95F;
		end
		32'h00001588: begin
				q			<=			16'h18B7;
		end
		32'h0000158A: begin
				q			<=			16'h0001;
		end
		32'h0000158C: begin
				q			<=			16'h8893;
		end
		32'h0000158E: begin
				q			<=			16'hE1C8;
		end
		32'h00001590: begin
				q			<=			16'hF06F;
		end
		32'h00001592: begin
				q			<=			16'hF89F;
		end
		32'h00001594: begin
				q			<=			16'h0000;
		end
		32'h00001596: begin
				q			<=			16'h0000;
		end
		32'h00001598: begin
				q			<=			16'h0113;
		end
		32'h0000159A: begin
				q			<=			16'hFE01;
		end
		32'h0000159C: begin
				q			<=			16'h2E23;
		end
		32'h0000159E: begin
				q			<=			16'h0011;
		end
		32'h000015A0: begin
				q			<=			16'h2C23;
		end
		32'h000015A2: begin
				q			<=			16'h0081;
		end
		32'h000015A4: begin
				q			<=			16'h2A23;
		end
		32'h000015A6: begin
				q			<=			16'h0091;
		end
		32'h000015A8: begin
				q			<=			16'h2823;
		end
		32'h000015AA: begin
				q			<=			16'h0121;
		end
		32'h000015AC: begin
				q			<=			16'h2623;
		end
		32'h000015AE: begin
				q			<=			16'h0131;
		end
		32'h000015B0: begin
				q			<=			16'h0413;
		end
		32'h000015B2: begin
				q			<=			16'h0005;
		end
		32'h000015B4: begin
				q			<=			16'h8493;
		end
		32'h000015B6: begin
				q			<=			16'h0005;
		end
		32'h000015B8: begin
				q			<=			16'h0513;
		end
		32'h000015BA: begin
				q			<=			16'hFFC5;
		end
		32'h000015BC: begin
				q			<=			16'h0713;
		end
		32'h000015BE: begin
				q			<=			16'h0030;
		end
		32'h000015C0: begin
				q			<=			16'h0793;
		end
		32'h000015C2: begin
				q			<=			16'h0080;
		end
		32'h000015C4: begin
				q			<=			16'h7A63;
		end
		32'h000015C6: begin
				q			<=			16'h00B7;
		end
		32'h000015C8: begin
				q			<=			16'h07B3;
		end
		32'h000015CA: begin
				q			<=			16'h40B0;
		end
		32'h000015CC: begin
				q			<=			16'hF793;
		end
		32'h000015CE: begin
				q			<=			16'h0037;
		end
		32'h000015D0: begin
				q			<=			16'h8713;
		end
		32'h000015D2: begin
				q			<=			16'h0045;
		end
		32'h000015D4: begin
				q			<=			16'h87B3;
		end
		32'h000015D6: begin
				q			<=			16'h00E7;
		end
		32'h000015D8: begin
				q			<=			16'h0E63;
		end
		32'h000015DA: begin
				q			<=			16'h0204;
		end
		32'h000015DC: begin
				q			<=			16'h2703;
		end
		32'h000015DE: begin
				q			<=			16'hFFC4;
		end
		32'h000015E0: begin
				q			<=			16'h6263;
		end
		32'h000015E2: begin
				q			<=			16'h04F7;
		end
		32'h000015E4: begin
				q			<=			16'h0733;
		end
		32'h000015E6: begin
				q			<=			16'h40F7;
		end
		32'h000015E8: begin
				q			<=			16'h0693;
		end
		32'h000015EA: begin
				q			<=			16'h0070;
		end
		32'h000015EC: begin
				q			<=			16'h0993;
		end
		32'h000015EE: begin
				q			<=			16'h0004;
		end
		32'h000015F0: begin
				q			<=			16'hE663;
		end
		32'h000015F2: begin
				q			<=			16'h06E6;
		end
		32'h000015F4: begin
				q			<=			16'h8513;
		end
		32'h000015F6: begin
				q			<=			16'h0009;
		end
		32'h000015F8: begin
				q			<=			16'h2083;
		end
		32'h000015FA: begin
				q			<=			16'h01C1;
		end
		32'h000015FC: begin
				q			<=			16'h2403;
		end
		32'h000015FE: begin
				q			<=			16'h0181;
		end
		32'h00001600: begin
				q			<=			16'h2483;
		end
		32'h00001602: begin
				q			<=			16'h0141;
		end
		32'h00001604: begin
				q			<=			16'h2903;
		end
		32'h00001606: begin
				q			<=			16'h0101;
		end
		32'h00001608: begin
				q			<=			16'h2983;
		end
		32'h0000160A: begin
				q			<=			16'h00C1;
		end
		32'h0000160C: begin
				q			<=			16'h0113;
		end
		32'h0000160E: begin
				q			<=			16'h0201;
		end
		32'h00001610: begin
				q			<=			16'h8067;
		end
		32'h00001612: begin
				q			<=			16'h0000;
		end
		32'h00001614: begin
				q			<=			16'h8513;
		end
		32'h00001616: begin
				q			<=			16'h0004;
		end
		32'h00001618: begin
				q			<=			16'hF0EF;
		end
		32'h0000161A: begin
				q			<=			16'hD91F;
		end
		32'h0000161C: begin
				q			<=			16'h0993;
		end
		32'h0000161E: begin
				q			<=			16'h0005;
		end
		32'h00001620: begin
				q			<=			16'hF06F;
		end
		32'h00001622: begin
				q			<=			16'hFD5F;
		end
		32'h00001624: begin
				q			<=			16'h0913;
		end
		32'h00001626: begin
				q			<=			16'hFFC7;
		end
		32'h00001628: begin
				q			<=			16'h8513;
		end
		32'h0000162A: begin
				q			<=			16'h0004;
		end
		32'h0000162C: begin
				q			<=			16'hF0EF;
		end
		32'h0000162E: begin
				q			<=			16'hD7DF;
		end
		32'h00001630: begin
				q			<=			16'h0993;
		end
		32'h00001632: begin
				q			<=			16'h0005;
		end
		32'h00001634: begin
				q			<=			16'h00E3;
		end
		32'h00001636: begin
				q			<=			16'hFC05;
		end
		32'h00001638: begin
				q			<=			16'h8613;
		end
		32'h0000163A: begin
				q			<=			16'h0004;
		end
		32'h0000163C: begin
				q			<=			16'h7463;
		end
		32'h0000163E: begin
				q			<=			16'h0099;
		end
		32'h00001640: begin
				q			<=			16'h0613;
		end
		32'h00001642: begin
				q			<=			16'h0009;
		end
		32'h00001644: begin
				q			<=			16'h0593;
		end
		32'h00001646: begin
				q			<=			16'h0004;
		end
		32'h00001648: begin
				q			<=			16'h8513;
		end
		32'h0000164A: begin
				q			<=			16'h0009;
		end
		32'h0000164C: begin
				q			<=			16'h10EF;
		end
		32'h0000164E: begin
				q			<=			16'h4AC0;
		end
		32'h00001650: begin
				q			<=			16'h0513;
		end
		32'h00001652: begin
				q			<=			16'h0004;
		end
		32'h00001654: begin
				q			<=			16'hF0EF;
		end
		32'h00001656: begin
				q			<=			16'hE75F;
		end
		32'h00001658: begin
				q			<=			16'hF06F;
		end
		32'h0000165A: begin
				q			<=			16'hF9DF;
		end
		32'h0000165C: begin
				q			<=			16'h0533;
		end
		32'h0000165E: begin
				q			<=			16'h00F5;
		end
		32'h00001660: begin
				q			<=			16'h2E23;
		end
		32'h00001662: begin
				q			<=			16'hFEF4;
		end
		32'h00001664: begin
				q			<=			16'h2023;
		end
		32'h00001666: begin
				q			<=			16'h00E5;
		end
		32'h00001668: begin
				q			<=			16'h0513;
		end
		32'h0000166A: begin
				q			<=			16'h0045;
		end
		32'h0000166C: begin
				q			<=			16'hF0EF;
		end
		32'h0000166E: begin
				q			<=			16'hE5DF;
		end
		32'h00001670: begin
				q			<=			16'hF06F;
		end
		32'h00001672: begin
				q			<=			16'hF85F;
		end
		32'h00001674: begin
				q			<=			16'h0000;
		end
		32'h00001676: begin
				q			<=			16'h0000;
		end
		32'h00001678: begin
				q			<=			16'h0113;
		end
		32'h0000167A: begin
				q			<=			16'hFF01;
		end
		32'h0000167C: begin
				q			<=			16'h2623;
		end
		32'h0000167E: begin
				q			<=			16'h0011;
		end
		32'h00001680: begin
				q			<=			16'h2423;
		end
		32'h00001682: begin
				q			<=			16'h0081;
		end
		32'h00001684: begin
				q			<=			16'h2223;
		end
		32'h00001686: begin
				q			<=			16'h0091;
		end
		32'h00001688: begin
				q			<=			16'h04B3;
		end
		32'h0000168A: begin
				q			<=			16'h02B5;
		end
		32'h0000168C: begin
				q			<=			16'h8513;
		end
		32'h0000168E: begin
				q			<=			16'h0004;
		end
		32'h00001690: begin
				q			<=			16'hF0EF;
		end
		32'h00001692: begin
				q			<=			16'hD19F;
		end
		32'h00001694: begin
				q			<=			16'h0413;
		end
		32'h00001696: begin
				q			<=			16'h0005;
		end
		32'h00001698: begin
				q			<=			16'h0A63;
		end
		32'h0000169A: begin
				q			<=			16'h0005;
		end
		32'h0000169C: begin
				q			<=			16'h8613;
		end
		32'h0000169E: begin
				q			<=			16'h0004;
		end
		32'h000016A0: begin
				q			<=			16'h0593;
		end
		32'h000016A2: begin
				q			<=			16'h0000;
		end
		32'h000016A4: begin
				q			<=			16'h1097;
		end
		32'h000016A6: begin
				q			<=			16'h0000;
		end
		32'h000016A8: begin
				q			<=			16'h80E7;
		end
		32'h000016AA: begin
				q			<=			16'h5400;
		end
		32'h000016AC: begin
				q			<=			16'h0513;
		end
		32'h000016AE: begin
				q			<=			16'h0004;
		end
		32'h000016B0: begin
				q			<=			16'h2083;
		end
		32'h000016B2: begin
				q			<=			16'h00C1;
		end
		32'h000016B4: begin
				q			<=			16'h2403;
		end
		32'h000016B6: begin
				q			<=			16'h0081;
		end
		32'h000016B8: begin
				q			<=			16'h2483;
		end
		32'h000016BA: begin
				q			<=			16'h0041;
		end
		32'h000016BC: begin
				q			<=			16'h0113;
		end
		32'h000016BE: begin
				q			<=			16'h0101;
		end
		32'h000016C0: begin
				q			<=			16'h8067;
		end
		32'h000016C2: begin
				q			<=			16'h0000;
		end
		32'h000016C4: begin
				q			<=			16'h0000;
		end
		32'h000016C6: begin
				q			<=			16'h0000;
		end
		32'h000016C8: begin
				q			<=			16'h0113;
		end
		32'h000016CA: begin
				q			<=			16'hFF01;
		end
		32'h000016CC: begin
				q			<=			16'h2623;
		end
		32'h000016CE: begin
				q			<=			16'h0011;
		end
		32'h000016D0: begin
				q			<=			16'hF0EF;
		end
		32'h000016D2: begin
				q			<=			16'hDF9F;
		end
		32'h000016D4: begin
				q			<=			16'h2083;
		end
		32'h000016D6: begin
				q			<=			16'h00C1;
		end
		32'h000016D8: begin
				q			<=			16'h0113;
		end
		32'h000016DA: begin
				q			<=			16'h0101;
		end
		32'h000016DC: begin
				q			<=			16'h8067;
		end
		32'h000016DE: begin
				q			<=			16'h0000;
		end
		32'h000016E0: begin
				q			<=			16'h0000;
		end
		32'h000016E2: begin
				q			<=			16'h0000;
		end
		32'h000016E4: begin
				q			<=			16'h0793;
		end
		32'h000016E6: begin
				q			<=			16'h0030;
		end
		32'h000016E8: begin
				q			<=			16'h0893;
		end
		32'h000016EA: begin
				q			<=			16'h0080;
		end
		32'h000016EC: begin
				q			<=			16'hFA63;
		end
		32'h000016EE: begin
				q			<=			16'h00B7;
		end
		32'h000016F0: begin
				q			<=			16'h08B3;
		end
		32'h000016F2: begin
				q			<=			16'h40B0;
		end
		32'h000016F4: begin
				q			<=			16'hF893;
		end
		32'h000016F6: begin
				q			<=			16'h0038;
		end
		32'h000016F8: begin
				q			<=			16'h8593;
		end
		32'h000016FA: begin
				q			<=			16'h0045;
		end
		32'h000016FC: begin
				q			<=			16'h88B3;
		end
		32'h000016FE: begin
				q			<=			16'h00B8;
		end
		32'h00001700: begin
				q			<=			16'h0813;
		end
		32'h00001702: begin
				q			<=			16'hFFF5;
		end
		32'h00001704: begin
				q			<=			16'h77B3;
		end
		32'h00001706: begin
				q			<=			16'h00A8;
		end
		32'h00001708: begin
				q			<=			16'h9663;
		end
		32'h0000170A: begin
				q			<=			16'h1807;
		end
		32'h0000170C: begin
				q			<=			16'h0863;
		end
		32'h0000170E: begin
				q			<=			16'h1805;
		end
		32'h00001710: begin
				q			<=			16'h0113;
		end
		32'h00001712: begin
				q			<=			16'hFF01;
		end
		32'h00001714: begin
				q			<=			16'h2623;
		end
		32'h00001716: begin
				q			<=			16'h0081;
		end
		32'h00001718: begin
				q			<=			16'h0413;
		end
		32'h0000171A: begin
				q			<=			16'h0101;
		end
		32'h0000171C: begin
				q			<=			16'h17B7;
		end
		32'h0000171E: begin
				q			<=			16'h0001;
		end
		32'h00001720: begin
				q			<=			16'h8593;
		end
		32'h00001722: begin
				q			<=			16'hE1C7;
		end
		32'h00001724: begin
				q			<=			16'h1337;
		end
		32'h00001726: begin
				q			<=			16'h0001;
		end
		32'h00001728: begin
				q			<=			16'h0E93;
		end
		32'h0000172A: begin
				q			<=			16'hFFC0;
		end
		32'h0000172C: begin
				q			<=			16'h0E13;
		end
		32'h0000172E: begin
				q			<=			16'hFE00;
		end
		32'h00001730: begin
				q			<=			16'h006F;
		end
		32'h00001732: begin
				q			<=			16'h1000;
		end
		32'h00001734: begin
				q			<=			16'h2603;
		end
		32'h00001736: begin
				q			<=			16'h8EC3;
		end
		32'h00001738: begin
				q			<=			16'h8733;
		end
		32'h0000173A: begin
				q			<=			16'h40CE;
		end
		32'h0000173C: begin
				q			<=			16'h7733;
		end
		32'h0000173E: begin
				q			<=			16'h0107;
		end
		32'h00001740: begin
				q			<=			16'h0733;
		end
		32'h00001742: begin
				q			<=			16'h0117;
		end
		32'h00001744: begin
				q			<=			16'h06B3;
		end
		32'h00001746: begin
				q			<=			16'h40CE;
		end
		32'h00001748: begin
				q			<=			16'h06B3;
		end
		32'h0000174A: begin
				q			<=			16'h00D4;
		end
		32'h0000174C: begin
				q			<=			16'hEC63;
		end
		32'h0000174E: begin
				q			<=			16'h14E6;
		end
		32'h00001750: begin
				q			<=			16'h07B3;
		end
		32'h00001752: begin
				q			<=			16'h00E6;
		end
		32'h00001754: begin
				q			<=			16'h2623;
		end
		32'h00001756: begin
				q			<=			16'h8EF3;
		end
		32'h00001758: begin
				q			<=			16'hA023;
		end
		32'h0000175A: begin
				q			<=			16'h00C5;
		end
		32'h0000175C: begin
				q			<=			16'h2023;
		end
		32'h0000175E: begin
				q			<=			16'h00E6;
		end
		32'h00001760: begin
				q			<=			16'h2223;
		end
		32'h00001762: begin
				q			<=			16'h0006;
		end
		32'h00001764: begin
				q			<=			16'h0513;
		end
		32'h00001766: begin
				q			<=			16'h0046;
		end
		32'h00001768: begin
				q			<=			16'h06B3;
		end
		32'h0000176A: begin
				q			<=			16'h40A0;
		end
		32'h0000176C: begin
				q			<=			16'hF7B3;
		end
		32'h0000176E: begin
				q			<=			16'h0106;
		end
		32'h00001770: begin
				q			<=			16'h9C63;
		end
		32'h00001772: begin
				q			<=			16'h0807;
		end
		32'h00001774: begin
				q			<=			16'h86B3;
		end
		32'h00001776: begin
				q			<=			16'h00F8;
		end
		32'h00001778: begin
				q			<=			16'h7463;
		end
		32'h0000177A: begin
				q			<=			16'h04D7;
		end
		32'h0000177C: begin
				q			<=			16'h2703;
		end
		32'h0000177E: begin
				q			<=			16'h0006;
		end
		32'h00001780: begin
				q			<=			16'h0733;
		end
		32'h00001782: begin
				q			<=			16'h00E6;
		end
		32'h00001784: begin
				q			<=			16'h2F83;
		end
		32'h00001786: begin
				q			<=			16'h8EC3;
		end
		32'h00001788: begin
				q			<=			16'h9063;
		end
		32'h0000178A: begin
				q			<=			16'h0AEF;
		end
		32'h0000178C: begin
				q			<=			16'h1737;
		end
		32'h0000178E: begin
				q			<=			16'h0001;
		end
		32'h00001790: begin
				q			<=			16'h2703;
		end
		32'h00001792: begin
				q			<=			16'h8EC7;
		end
		32'h00001794: begin
				q			<=			16'h0733;
		end
		32'h00001796: begin
				q			<=			16'h40E4;
		end
		32'h00001798: begin
				q			<=			16'h0713;
		end
		32'h0000179A: begin
				q			<=			16'hFE07;
		end
		32'h0000179C: begin
				q			<=			16'h2803;
		end
		32'h0000179E: begin
				q			<=			16'h0006;
		end
		32'h000017A0: begin
				q			<=			16'h8833;
		end
		32'h000017A2: begin
				q			<=			16'h4106;
		end
		32'h000017A4: begin
				q			<=			16'h6463;
		end
		32'h000017A6: begin
				q			<=			16'h1107;
		end
		32'h000017A8: begin
				q			<=			16'h0F33;
		end
		32'h000017AA: begin
				q			<=			16'h00F6;
		end
		32'h000017AC: begin
				q			<=			16'h0F33;
		end
		32'h000017AE: begin
				q			<=			16'h011F;
		end
		32'h000017B0: begin
				q			<=			16'h1737;
		end
		32'h000017B2: begin
				q			<=			16'h0001;
		end
		32'h000017B4: begin
				q			<=			16'h2623;
		end
		32'h000017B6: begin
				q			<=			16'h8FE7;
		end
		32'h000017B8: begin
				q			<=			16'h2023;
		end
		32'h000017BA: begin
				q			<=			16'h00D6;
		end
		32'h000017BC: begin
				q			<=			16'h8713;
		end
		32'h000017BE: begin
				q			<=			16'h0006;
		end
		32'h000017C0: begin
				q			<=			16'h8E63;
		end
		32'h000017C2: begin
				q			<=			16'h0807;
		end
		32'h000017C4: begin
				q			<=			16'h2023;
		end
		32'h000017C6: begin
				q			<=			16'h00F6;
		end
		32'h000017C8: begin
				q			<=			16'h06B3;
		end
		32'h000017CA: begin
				q			<=			16'h00F6;
		end
		32'h000017CC: begin
				q			<=			16'h8513;
		end
		32'h000017CE: begin
				q			<=			16'h0006;
		end
		32'h000017D0: begin
				q			<=			16'h07B3;
		end
		32'h000017D2: begin
				q			<=			16'h40F7;
		end
		32'h000017D4: begin
				q			<=			16'h8713;
		end
		32'h000017D6: begin
				q			<=			16'h0088;
		end
		32'h000017D8: begin
				q			<=			16'h7C63;
		end
		32'h000017DA: begin
				q			<=			16'h06F7;
		end
		32'h000017DC: begin
				q			<=			16'h86B3;
		end
		32'h000017DE: begin
				q			<=			16'h00D8;
		end
		32'h000017E0: begin
				q			<=			16'h87B3;
		end
		32'h000017E2: begin
				q			<=			16'h4117;
		end
		32'h000017E4: begin
				q			<=			16'hA023;
		end
		32'h000017E6: begin
				q			<=			16'h00F6;
		end
		32'h000017E8: begin
				q			<=			16'h2783;
		end
		32'h000017EA: begin
				q			<=			16'h0046;
		end
		32'h000017EC: begin
				q			<=			16'hA223;
		end
		32'h000017EE: begin
				q			<=			16'h00F6;
		end
		32'h000017F0: begin
				q			<=			16'h2223;
		end
		32'h000017F2: begin
				q			<=			16'h00D6;
		end
		32'h000017F4: begin
				q			<=			16'h2023;
		end
		32'h000017F6: begin
				q			<=			16'h0115;
		end
		32'h000017F8: begin
				q			<=			16'h0513;
		end
		32'h000017FA: begin
				q			<=			16'h0045;
		end
		32'h000017FC: begin
				q			<=			16'h2403;
		end
		32'h000017FE: begin
				q			<=			16'h00C1;
		end
		32'h00001800: begin
				q			<=			16'h0113;
		end
		32'h00001802: begin
				q			<=			16'h0101;
		end
		32'h00001804: begin
				q			<=			16'h8067;
		end
		32'h00001806: begin
				q			<=			16'h0000;
		end
		32'h00001808: begin
				q			<=			16'h0793;
		end
		32'h0000180A: begin
				q			<=			16'h00C6;
		end
		32'h0000180C: begin
				q			<=			16'h07B3;
		end
		32'h0000180E: begin
				q			<=			16'h40F0;
		end
		32'h00001810: begin
				q			<=			16'hF7B3;
		end
		32'h00001812: begin
				q			<=			16'h0107;
		end
		32'h00001814: begin
				q			<=			16'h8793;
		end
		32'h00001816: begin
				q			<=			16'h0087;
		end
		32'h00001818: begin
				q			<=			16'h2683;
		end
		32'h0000181A: begin
				q			<=			16'h0046;
		end
		32'h0000181C: begin
				q			<=			16'h8CE3;
		end
		32'h0000181E: begin
				q			<=			16'hF406;
		end
		32'h00001820: begin
				q			<=			16'h86B3;
		end
		32'h00001822: begin
				q			<=			16'h0117;
		end
		32'h00001824: begin
				q			<=			16'h7EE3;
		end
		32'h00001826: begin
				q			<=			16'hF8D7;
		end
		32'h00001828: begin
				q			<=			16'hA783;
		end
		32'h0000182A: begin
				q			<=			16'h0005;
		end
		32'h0000182C: begin
				q			<=			16'h8593;
		end
		32'h0000182E: begin
				q			<=			16'h0047;
		end
		32'h00001830: begin
				q			<=			16'hA603;
		end
		32'h00001832: begin
				q			<=			16'h0005;
		end
		32'h00001834: begin
				q			<=			16'h00E3;
		end
		32'h00001836: begin
				q			<=			16'hF006;
		end
		32'h00001838: begin
				q			<=			16'h2703;
		end
		32'h0000183A: begin
				q			<=			16'h0006;
		end
		32'h0000183C: begin
				q			<=			16'h0513;
		end
		32'h0000183E: begin
				q			<=			16'h0046;
		end
		32'h00001840: begin
				q			<=			16'h06B3;
		end
		32'h00001842: begin
				q			<=			16'h40A0;
		end
		32'h00001844: begin
				q			<=			16'hF7B3;
		end
		32'h00001846: begin
				q			<=			16'h0106;
		end
		32'h00001848: begin
				q			<=			16'h88E3;
		end
		32'h0000184A: begin
				q			<=			16'hFC07;
		end
		32'h0000184C: begin
				q			<=			16'hF06F;
		end
		32'h0000184E: begin
				q			<=			16'hFBDF;
		end
		32'h00001850: begin
				q			<=			16'hA023;
		end
		32'h00001852: begin
				q			<=			16'h00F6;
		end
		32'h00001854: begin
				q			<=			16'h8513;
		end
		32'h00001856: begin
				q			<=			16'h0046;
		end
		32'h00001858: begin
				q			<=			16'hF06F;
		end
		32'h0000185A: begin
				q			<=			16'hFA5F;
		end
		32'h0000185C: begin
				q			<=			16'h8793;
		end
		32'h0000185E: begin
				q			<=			16'h0088;
		end
		32'h00001860: begin
				q			<=			16'hF463;
		end
		32'h00001862: begin
				q			<=			16'h02E7;
		end
		32'h00001864: begin
				q			<=			16'h2683;
		end
		32'h00001866: begin
				q			<=			16'h0046;
		end
		32'h00001868: begin
				q			<=			16'h07B3;
		end
		32'h0000186A: begin
				q			<=			16'h0116;
		end
		32'h0000186C: begin
				q			<=			16'hA023;
		end
		32'h0000186E: begin
				q			<=			16'h00F5;
		end
		32'h00001870: begin
				q			<=			16'h0733;
		end
		32'h00001872: begin
				q			<=			16'h4117;
		end
		32'h00001874: begin
				q			<=			16'hA023;
		end
		32'h00001876: begin
				q			<=			16'h00E7;
		end
		32'h00001878: begin
				q			<=			16'hA783;
		end
		32'h0000187A: begin
				q			<=			16'h0005;
		end
		32'h0000187C: begin
				q			<=			16'hA223;
		end
		32'h0000187E: begin
				q			<=			16'h00D7;
		end
		32'h00001880: begin
				q			<=			16'h0513;
		end
		32'h00001882: begin
				q			<=			16'h0006;
		end
		32'h00001884: begin
				q			<=			16'hF06F;
		end
		32'h00001886: begin
				q			<=			16'hF71F;
		end
		32'h00001888: begin
				q			<=			16'h2783;
		end
		32'h0000188A: begin
				q			<=			16'h0046;
		end
		32'h0000188C: begin
				q			<=			16'hA023;
		end
		32'h0000188E: begin
				q			<=			16'h00F5;
		end
		32'h00001890: begin
				q			<=			16'hF06F;
		end
		32'h00001892: begin
				q			<=			16'hF6DF;
		end
		32'h00001894: begin
				q			<=			16'h0513;
		end
		32'h00001896: begin
				q			<=			16'h0000;
		end
		32'h00001898: begin
				q			<=			16'h8067;
		end
		32'h0000189A: begin
				q			<=			16'h0000;
		end
		32'h0000189C: begin
				q			<=			16'h0513;
		end
		32'h0000189E: begin
				q			<=			16'h0000;
		end
		32'h000018A0: begin
				q			<=			16'h8067;
		end
		32'h000018A2: begin
				q			<=			16'h0000;
		end
		32'h000018A4: begin
				q			<=			16'h0513;
		end
		32'h000018A6: begin
				q			<=			16'h0000;
		end
		32'h000018A8: begin
				q			<=			16'hF06F;
		end
		32'h000018AA: begin
				q			<=			16'hF55F;
		end
		32'h000018AC: begin
				q			<=			16'h0513;
		end
		32'h000018AE: begin
				q			<=			16'h0000;
		end
		32'h000018B0: begin
				q			<=			16'hF06F;
		end
		32'h000018B2: begin
				q			<=			16'hF4DF;
		end
		32'h000018B4: begin
				q			<=			16'h0000;
		end
		32'h000018B6: begin
				q			<=			16'h0000;
		end
		32'h000018B8: begin
				q			<=			16'h0113;
		end
		32'h000018BA: begin
				q			<=			16'hFF01;
		end
		32'h000018BC: begin
				q			<=			16'h2623;
		end
		32'h000018BE: begin
				q			<=			16'h0011;
		end
		32'h000018C0: begin
				q			<=			16'h0593;
		end
		32'h000018C2: begin
				q			<=			16'h0005;
		end
		32'h000018C4: begin
				q			<=			16'h0513;
		end
		32'h000018C6: begin
				q			<=			16'h0800;
		end
		32'h000018C8: begin
				q			<=			16'hF0EF;
		end
		32'h000018CA: begin
				q			<=			16'hE1DF;
		end
		32'h000018CC: begin
				q			<=			16'h2083;
		end
		32'h000018CE: begin
				q			<=			16'h00C1;
		end
		32'h000018D0: begin
				q			<=			16'h0113;
		end
		32'h000018D2: begin
				q			<=			16'h0101;
		end
		32'h000018D4: begin
				q			<=			16'h8067;
		end
		32'h000018D6: begin
				q			<=			16'h0000;
		end
		32'h000018D8: begin
				q			<=			16'h0000;
		end
		32'h000018DA: begin
				q			<=			16'h0000;
		end
		32'h000018DC: begin
				q			<=			16'h0113;
		end
		32'h000018DE: begin
				q			<=			16'hFF01;
		end
		32'h000018E0: begin
				q			<=			16'h2623;
		end
		32'h000018E2: begin
				q			<=			16'h0011;
		end
		32'h000018E4: begin
				q			<=			16'h07B3;
		end
		32'h000018E6: begin
				q			<=			16'h40A0;
		end
		32'h000018E8: begin
				q			<=			16'hF793;
		end
		32'h000018EA: begin
				q			<=			16'h07F7;
		end
		32'h000018EC: begin
				q			<=			16'h85B3;
		end
		32'h000018EE: begin
				q			<=			16'h00A7;
		end
		32'h000018F0: begin
				q			<=			16'h0513;
		end
		32'h000018F2: begin
				q			<=			16'h0800;
		end
		32'h000018F4: begin
				q			<=			16'hF0EF;
		end
		32'h000018F6: begin
				q			<=			16'hDF1F;
		end
		32'h000018F8: begin
				q			<=			16'h2083;
		end
		32'h000018FA: begin
				q			<=			16'h00C1;
		end
		32'h000018FC: begin
				q			<=			16'h0113;
		end
		32'h000018FE: begin
				q			<=			16'h0101;
		end
		32'h00001900: begin
				q			<=			16'h8067;
		end
		32'h00001902: begin
				q			<=			16'h0000;
		end
		32'h00001904: begin
				q			<=			16'h0000;
		end
		32'h00001906: begin
				q			<=			16'h0000;
		end
		32'h00001908: begin
				q			<=			16'h0113;
		end
		32'h0000190A: begin
				q			<=			16'hFC01;
		end
		32'h0000190C: begin
				q			<=			16'h2E23;
		end
		32'h0000190E: begin
				q			<=			16'h0211;
		end
		32'h00001910: begin
				q			<=			16'h2C23;
		end
		32'h00001912: begin
				q			<=			16'h0281;
		end
		32'h00001914: begin
				q			<=			16'h0413;
		end
		32'h00001916: begin
				q			<=			16'h0005;
		end
		32'h00001918: begin
				q			<=			16'h0613;
		end
		32'h0000191A: begin
				q			<=			16'h0280;
		end
		32'h0000191C: begin
				q			<=			16'h0593;
		end
		32'h0000191E: begin
				q			<=			16'h0000;
		end
		32'h00001920: begin
				q			<=			16'h0513;
		end
		32'h00001922: begin
				q			<=			16'h0081;
		end
		32'h00001924: begin
				q			<=			16'h1097;
		end
		32'h00001926: begin
				q			<=			16'h0000;
		end
		32'h00001928: begin
				q			<=			16'h80E7;
		end
		32'h0000192A: begin
				q			<=			16'h2C00;
		end
		32'h0000192C: begin
				q			<=			16'h17B7;
		end
		32'h0000192E: begin
				q			<=			16'h0001;
		end
		32'h00001930: begin
				q			<=			16'hA783;
		end
		32'h00001932: begin
				q			<=			16'hE1C7;
		end
		32'h00001934: begin
				q			<=			16'h8863;
		end
		32'h00001936: begin
				q			<=			16'h0807;
		end
		32'h00001938: begin
				q			<=			16'h1737;
		end
		32'h0000193A: begin
				q			<=			16'h0001;
		end
		32'h0000193C: begin
				q			<=			16'h2503;
		end
		32'h0000193E: begin
				q			<=			16'h8EC7;
		end
		32'h00001940: begin
				q			<=			16'h0593;
		end
		32'h00001942: begin
				q			<=			16'h0000;
		end
		32'h00001944: begin
				q			<=			16'h0693;
		end
		32'h00001946: begin
				q			<=			16'h0000;
		end
		32'h00001948: begin
				q			<=			16'h006F;
		end
		32'h0000194A: begin
				q			<=			16'h0140;
		end
		32'h0000194C: begin
				q			<=			16'h2623;
		end
		32'h0000194E: begin
				q			<=			16'h02C1;
		end
		32'h00001950: begin
				q			<=			16'hA703;
		end
		32'h00001952: begin
				q			<=			16'h0047;
		end
		32'h00001954: begin
				q			<=			16'h0263;
		end
		32'h00001956: begin
				q			<=			16'h0207;
		end
		32'h00001958: begin
				q			<=			16'h0793;
		end
		32'h0000195A: begin
				q			<=			16'h0007;
		end
		32'h0000195C: begin
				q			<=			16'hA603;
		end
		32'h0000195E: begin
				q			<=			16'h0007;
		end
		32'h00001960: begin
				q			<=			16'h86B3;
		end
		32'h00001962: begin
				q			<=			16'h00C6;
		end
		32'h00001964: begin
				q			<=			16'h8593;
		end
		32'h00001966: begin
				q			<=			16'h0015;
		end
		32'h00001968: begin
				q			<=			16'hA703;
		end
		32'h0000196A: begin
				q			<=			16'h0047;
		end
		32'h0000196C: begin
				q			<=			16'h16E3;
		end
		32'h0000196E: begin
				q			<=			16'hFE07;
		end
		32'h00001970: begin
				q			<=			16'h8733;
		end
		32'h00001972: begin
				q			<=			16'h00C7;
		end
		32'h00001974: begin
				q			<=			16'h0CE3;
		end
		32'h00001976: begin
				q			<=			16'hFCE5;
		end
		32'h00001978: begin
				q			<=			16'h17B7;
		end
		32'h0000197A: begin
				q			<=			16'h0001;
		end
		32'h0000197C: begin
				q			<=			16'hA783;
		end
		32'h0000197E: begin
				q			<=			16'h8EC7;
		end
		32'h00001980: begin
				q			<=			16'h0737;
		end
		32'h00001982: begin
				q			<=			16'h0100;
		end
		32'h00001984: begin
				q			<=			16'h0713;
		end
		32'h00001986: begin
				q			<=			16'h0007;
		end
		32'h00001988: begin
				q			<=			16'h87B3;
		end
		32'h0000198A: begin
				q			<=			16'h40E7;
		end
		32'h0000198C: begin
				q			<=			16'h2423;
		end
		32'h0000198E: begin
				q			<=			16'h00F1;
		end
		32'h00001990: begin
				q			<=			16'h2423;
		end
		32'h00001992: begin
				q			<=			16'h02D1;
		end
		32'h00001994: begin
				q			<=			16'h86B3;
		end
		32'h00001996: begin
				q			<=			16'h40D7;
		end
		32'h00001998: begin
				q			<=			16'h2223;
		end
		32'h0000199A: begin
				q			<=			16'h02D1;
		end
		32'h0000199C: begin
				q			<=			16'h2623;
		end
		32'h0000199E: begin
				q			<=			16'h00B1;
		end
		32'h000019A0: begin
				q			<=			16'h0613;
		end
		32'h000019A2: begin
				q			<=			16'h0280;
		end
		32'h000019A4: begin
				q			<=			16'h0593;
		end
		32'h000019A6: begin
				q			<=			16'h0081;
		end
		32'h000019A8: begin
				q			<=			16'h0513;
		end
		32'h000019AA: begin
				q			<=			16'h0004;
		end
		32'h000019AC: begin
				q			<=			16'h10EF;
		end
		32'h000019AE: begin
				q			<=			16'h14C0;
		end
		32'h000019B0: begin
				q			<=			16'h0513;
		end
		32'h000019B2: begin
				q			<=			16'h0004;
		end
		32'h000019B4: begin
				q			<=			16'h2083;
		end
		32'h000019B6: begin
				q			<=			16'h03C1;
		end
		32'h000019B8: begin
				q			<=			16'h2403;
		end
		32'h000019BA: begin
				q			<=			16'h0381;
		end
		32'h000019BC: begin
				q			<=			16'h0113;
		end
		32'h000019BE: begin
				q			<=			16'h0401;
		end
		32'h000019C0: begin
				q			<=			16'h8067;
		end
		32'h000019C2: begin
				q			<=			16'h0000;
		end
		32'h000019C4: begin
				q			<=			16'h0593;
		end
		32'h000019C6: begin
				q			<=			16'h0000;
		end
		32'h000019C8: begin
				q			<=			16'h0693;
		end
		32'h000019CA: begin
				q			<=			16'h0000;
		end
		32'h000019CC: begin
				q			<=			16'hF06F;
		end
		32'h000019CE: begin
				q			<=			16'hFADF;
		end
		32'h000019D0: begin
				q			<=			16'h0000;
		end
		32'h000019D2: begin
				q			<=			16'h0000;
		end
		32'h000019D4: begin
				q			<=			16'h2503;
		end
		32'h000019D6: begin
				q			<=			16'hFFC5;
		end
		32'h000019D8: begin
				q			<=			16'h0513;
		end
		32'h000019DA: begin
				q			<=			16'hFFC5;
		end
		32'h000019DC: begin
				q			<=			16'h8067;
		end
		32'h000019DE: begin
				q			<=			16'h0000;
		end
		32'h000019E0: begin
				q			<=			16'h0000;
		end
		32'h000019E2: begin
				q			<=			16'h0000;
		end
		32'h000019E4: begin
				q			<=			16'h0513;
		end
		32'h000019E6: begin
				q			<=			16'h0000;
		end
		32'h000019E8: begin
				q			<=			16'h8067;
		end
		32'h000019EA: begin
				q			<=			16'h0000;
		end
		32'h000019EC: begin
				q			<=			16'h0000;
		end
		32'h000019EE: begin
				q			<=			16'h0000;
		end
		32'h000019F0: begin
				q			<=			16'h0113;
		end
		32'h000019F2: begin
				q			<=			16'hFD01;
		end
		32'h000019F4: begin
				q			<=			16'h2623;
		end
		32'h000019F6: begin
				q			<=			16'h0211;
		end
		32'h000019F8: begin
				q			<=			16'h2423;
		end
		32'h000019FA: begin
				q			<=			16'h0281;
		end
		32'h000019FC: begin
				q			<=			16'h0613;
		end
		32'h000019FE: begin
				q			<=			16'h1000;
		end
		32'h00001A00: begin
				q			<=			16'h0593;
		end
		32'h00001A02: begin
				q			<=			16'h0000;
		end
		32'h00001A04: begin
				q			<=			16'h1437;
		end
		32'h00001A06: begin
				q			<=			16'h0001;
		end
		32'h00001A08: begin
				q			<=			16'h0513;
		end
		32'h00001A0A: begin
				q			<=			16'hE3C4;
		end
		32'h00001A0C: begin
				q			<=			16'h1097;
		end
		32'h00001A0E: begin
				q			<=			16'h0000;
		end
		32'h00001A10: begin
				q			<=			16'h80E7;
		end
		32'h00001A12: begin
				q			<=			16'h1D80;
		end
		32'h00001A14: begin
				q			<=			16'h0793;
		end
		32'h00001A16: begin
				q			<=			16'h02F0;
		end
		32'h00001A18: begin
				q			<=			16'h0E23;
		end
		32'h00001A1A: begin
				q			<=			16'hE2F4;
		end
		32'h00001A1C: begin
				q			<=			16'h1537;
		end
		32'h00001A1E: begin
				q			<=			16'h0001;
		end
		32'h00001A20: begin
				q			<=			16'h0513;
		end
		32'h00001A22: begin
				q			<=			16'hF405;
		end
		32'h00001A24: begin
				q			<=			16'h00EF;
		end
		32'h00001A26: begin
				q			<=			16'h0910;
		end
		32'h00001A28: begin
				q			<=			16'h0793;
		end
		32'h00001A2A: begin
				q			<=			16'h0005;
		end
		32'h00001A2C: begin
				q			<=			16'h1737;
		end
		32'h00001A2E: begin
				q			<=			16'h0001;
		end
		32'h00001A30: begin
				q			<=			16'h2023;
		end
		32'h00001A32: begin
				q			<=			16'hE2A7;
		end
		32'h00001A34: begin
				q			<=			16'h0513;
		end
		32'h00001A36: begin
				q			<=			16'h0000;
		end
		32'h00001A38: begin
				q			<=			16'h8A63;
		end
		32'h00001A3A: begin
				q			<=			16'h0007;
		end
		32'h00001A3C: begin
				q			<=			16'h2083;
		end
		32'h00001A3E: begin
				q			<=			16'h02C1;
		end
		32'h00001A40: begin
				q			<=			16'h2403;
		end
		32'h00001A42: begin
				q			<=			16'h0281;
		end
		32'h00001A44: begin
				q			<=			16'h0113;
		end
		32'h00001A46: begin
				q			<=			16'h0301;
		end
		32'h00001A48: begin
				q			<=			16'h8067;
		end
		32'h00001A4A: begin
				q			<=			16'h0000;
		end
		32'h00001A4C: begin
				q			<=			16'h0593;
		end
		32'h00001A4E: begin
				q			<=			16'hE3C4;
		end
		32'h00001A50: begin
				q			<=			16'h0513;
		end
		32'h00001A52: begin
				q			<=			16'h00C1;
		end
		32'h00001A54: begin
				q			<=			16'h00EF;
		end
		32'h00001A56: begin
				q			<=			16'h48D0;
		end
		32'h00001A58: begin
				q			<=			16'h17B7;
		end
		32'h00001A5A: begin
				q			<=			16'h0001;
		end
		32'h00001A5C: begin
				q			<=			16'hA023;
		end
		32'h00001A5E: begin
				q			<=			16'hE2A7;
		end
		32'h00001A60: begin
				q			<=			16'h3513;
		end
		32'h00001A62: begin
				q			<=			16'h0015;
		end
		32'h00001A64: begin
				q			<=			16'hF06F;
		end
		32'h00001A66: begin
				q			<=			16'hFD9F;
		end
		32'h00001A68: begin
				q			<=			16'h0000;
		end
		32'h00001A6A: begin
				q			<=			16'h0000;
		end
		32'h00001A6C: begin
				q			<=			16'h0113;
		end
		32'h00001A6E: begin
				q			<=			16'hFD01;
		end
		32'h00001A70: begin
				q			<=			16'h2623;
		end
		32'h00001A72: begin
				q			<=			16'h0211;
		end
		32'h00001A74: begin
				q			<=			16'h2423;
		end
		32'h00001A76: begin
				q			<=			16'h0281;
		end
		32'h00001A78: begin
				q			<=			16'h2223;
		end
		32'h00001A7A: begin
				q			<=			16'h0291;
		end
		32'h00001A7C: begin
				q			<=			16'h0413;
		end
		32'h00001A7E: begin
				q			<=			16'h0005;
		end
		32'h00001A80: begin
				q			<=			16'h0593;
		end
		32'h00001A82: begin
				q			<=			16'h0005;
		end
		32'h00001A84: begin
				q			<=			16'h0513;
		end
		32'h00001A86: begin
				q			<=			16'h00C1;
		end
		32'h00001A88: begin
				q			<=			16'h00EF;
		end
		32'h00001A8A: begin
				q			<=			16'h4590;
		end
		32'h00001A8C: begin
				q			<=			16'h17B7;
		end
		32'h00001A8E: begin
				q			<=			16'h0001;
		end
		32'h00001A90: begin
				q			<=			16'hA023;
		end
		32'h00001A92: begin
				q			<=			16'hE2A7;
		end
		32'h00001A94: begin
				q			<=			16'h0863;
		end
		32'h00001A96: begin
				q			<=			16'h0205;
		end
		32'h00001A98: begin
				q			<=			16'h17B7;
		end
		32'h00001A9A: begin
				q			<=			16'h0001;
		end
		32'h00001A9C: begin
				q			<=			16'h0713;
		end
		32'h00001A9E: begin
				q			<=			16'h02F0;
		end
		32'h00001AA0: begin
				q			<=			16'h8E23;
		end
		32'h00001AA2: begin
				q			<=			16'hE2E7;
		end
		32'h00001AA4: begin
				q			<=			16'h8793;
		end
		32'h00001AA6: begin
				q			<=			16'hE3C7;
		end
		32'h00001AA8: begin
				q			<=			16'h80A3;
		end
		32'h00001AAA: begin
				q			<=			16'h0007;
		end
		32'h00001AAC: begin
				q			<=			16'h0513;
		end
		32'h00001AAE: begin
				q			<=			16'h0000;
		end
		32'h00001AB0: begin
				q			<=			16'h2083;
		end
		32'h00001AB2: begin
				q			<=			16'h02C1;
		end
		32'h00001AB4: begin
				q			<=			16'h2403;
		end
		32'h00001AB6: begin
				q			<=			16'h0281;
		end
		32'h00001AB8: begin
				q			<=			16'h2483;
		end
		32'h00001ABA: begin
				q			<=			16'h0241;
		end
		32'h00001ABC: begin
				q			<=			16'h0113;
		end
		32'h00001ABE: begin
				q			<=			16'h0301;
		end
		32'h00001AC0: begin
				q			<=			16'h8067;
		end
		32'h00001AC2: begin
				q			<=			16'h0000;
		end
		32'h00001AC4: begin
				q			<=			16'h0613;
		end
		32'h00001AC6: begin
				q			<=			16'h1000;
		end
		32'h00001AC8: begin
				q			<=			16'h0593;
		end
		32'h00001ACA: begin
				q			<=			16'h0000;
		end
		32'h00001ACC: begin
				q			<=			16'h14B7;
		end
		32'h00001ACE: begin
				q			<=			16'h0001;
		end
		32'h00001AD0: begin
				q			<=			16'h8513;
		end
		32'h00001AD2: begin
				q			<=			16'hE3C4;
		end
		32'h00001AD4: begin
				q			<=			16'h1097;
		end
		32'h00001AD6: begin
				q			<=			16'h0000;
		end
		32'h00001AD8: begin
				q			<=			16'h80E7;
		end
		32'h00001ADA: begin
				q			<=			16'h1100;
		end
		32'h00001ADC: begin
				q			<=			16'h0513;
		end
		32'h00001ADE: begin
				q			<=			16'h0004;
		end
		32'h00001AE0: begin
				q			<=			16'h10EF;
		end
		32'h00001AE2: begin
				q			<=			16'h34C0;
		end
		32'h00001AE4: begin
				q			<=			16'h0613;
		end
		32'h00001AE6: begin
				q			<=			16'h0005;
		end
		32'h00001AE8: begin
				q			<=			16'h0593;
		end
		32'h00001AEA: begin
				q			<=			16'h0004;
		end
		32'h00001AEC: begin
				q			<=			16'h8513;
		end
		32'h00001AEE: begin
				q			<=			16'hE3C4;
		end
		32'h00001AF0: begin
				q			<=			16'h10EF;
		end
		32'h00001AF2: begin
				q			<=			16'h39C0;
		end
		32'h00001AF4: begin
				q			<=			16'h0513;
		end
		32'h00001AF6: begin
				q			<=			16'h0010;
		end
		32'h00001AF8: begin
				q			<=			16'hF06F;
		end
		32'h00001AFA: begin
				q			<=			16'hFB9F;
		end
		32'h00001AFC: begin
				q			<=			16'h0000;
		end
		32'h00001AFE: begin
				q			<=			16'h0000;
		end
		32'h00001B00: begin
				q			<=			16'h0113;
		end
		32'h00001B02: begin
				q			<=			16'hFC01;
		end
		32'h00001B04: begin
				q			<=			16'h2E23;
		end
		32'h00001B06: begin
				q			<=			16'h0211;
		end
		32'h00001B08: begin
				q			<=			16'h2C23;
		end
		32'h00001B0A: begin
				q			<=			16'h0281;
		end
		32'h00001B0C: begin
				q			<=			16'h2A23;
		end
		32'h00001B0E: begin
				q			<=			16'h0291;
		end
		32'h00001B10: begin
				q			<=			16'h2823;
		end
		32'h00001B12: begin
				q			<=			16'h0321;
		end
		32'h00001B14: begin
				q			<=			16'h2623;
		end
		32'h00001B16: begin
				q			<=			16'h0331;
		end
		32'h00001B18: begin
				q			<=			16'h2423;
		end
		32'h00001B1A: begin
				q			<=			16'h0341;
		end
		32'h00001B1C: begin
				q			<=			16'h2223;
		end
		32'h00001B1E: begin
				q			<=			16'h0351;
		end
		32'h00001B20: begin
				q			<=			16'h2023;
		end
		32'h00001B22: begin
				q			<=			16'h0361;
		end
		32'h00001B24: begin
				q			<=			16'h15B7;
		end
		32'h00001B26: begin
				q			<=			16'h0001;
		end
		32'h00001B28: begin
				q			<=			16'h8593;
		end
		32'h00001B2A: begin
				q			<=			16'hE3C5;
		end
		32'h00001B2C: begin
				q			<=			16'h0513;
		end
		32'h00001B2E: begin
				q			<=			16'h00C1;
		end
		32'h00001B30: begin
				q			<=			16'h00EF;
		end
		32'h00001B32: begin
				q			<=			16'h3B10;
		end
		32'h00001B34: begin
				q			<=			16'h17B7;
		end
		32'h00001B36: begin
				q			<=			16'h0001;
		end
		32'h00001B38: begin
				q			<=			16'hA023;
		end
		32'h00001B3A: begin
				q			<=			16'hE2A7;
		end
		32'h00001B3C: begin
				q			<=			16'h1463;
		end
		32'h00001B3E: begin
				q			<=			16'h0A05;
		end
		32'h00001B40: begin
				q			<=			16'h0493;
		end
		32'h00001B42: begin
				q			<=			16'h03C0;
		end
		32'h00001B44: begin
				q			<=			16'h1437;
		end
		32'h00001B46: begin
				q			<=			16'h0001;
		end
		32'h00001B48: begin
				q			<=			16'h8993;
		end
		32'h00001B4A: begin
				q			<=			16'h0007;
		end
		32'h00001B4C: begin
				q			<=			16'h1A37;
		end
		32'h00001B4E: begin
				q			<=			16'h0001;
		end
		32'h00001B50: begin
				q			<=			16'h0B37;
		end
		32'h00001B52: begin
				q			<=			16'h0001;
		end
		32'h00001B54: begin
				q			<=			16'h1937;
		end
		32'h00001B56: begin
				q			<=			16'h0001;
		end
		32'h00001B58: begin
				q			<=			16'h0AB7;
		end
		32'h00001B5A: begin
				q			<=			16'h0001;
		end
		32'h00001B5C: begin
				q			<=			16'h006F;
		end
		32'h00001B5E: begin
				q			<=			16'h0300;
		end
		32'h00001B60: begin
				q			<=			16'h0693;
		end
		32'h00001B62: begin
				q			<=			16'hE2DA;
		end
		32'h00001B64: begin
				q			<=			16'h0613;
		end
		32'h00001B66: begin
				q			<=			16'hD68B;
		end
		32'h00001B68: begin
				q			<=			16'h0593;
		end
		32'h00001B6A: begin
				q			<=			16'h1000;
		end
		32'h00001B6C: begin
				q			<=			16'h0513;
		end
		32'h00001B6E: begin
				q			<=			16'hD1C9;
		end
		32'h00001B70: begin
				q			<=			16'h1097;
		end
		32'h00001B72: begin
				q			<=			16'h0000;
		end
		32'h00001B74: begin
				q			<=			16'h80E7;
		end
		32'h00001B76: begin
				q			<=			16'h1FC0;
		end
		32'h00001B78: begin
				q			<=			16'h0593;
		end
		32'h00001B7A: begin
				q			<=			16'h0010;
		end
		32'h00001B7C: begin
				q			<=			16'h0513;
		end
		32'h00001B7E: begin
				q			<=			16'hD1C9;
		end
		32'h00001B80: begin
				q			<=			16'hF0EF;
		end
		32'h00001B82: begin
				q			<=			16'h818F;
		end
		32'h00001B84: begin
				q			<=			16'h8493;
		end
		32'h00001B86: begin
				q			<=			16'hFFF4;
		end
		32'h00001B88: begin
				q			<=			16'h8E63;
		end
		32'h00001B8A: begin
				q			<=			16'h0404;
		end
		32'h00001B8C: begin
				q			<=			16'h0593;
		end
		32'h00001B8E: begin
				q			<=			16'hE244;
		end
		32'h00001B90: begin
				q			<=			16'h0513;
		end
		32'h00001B92: begin
				q			<=			16'h00C1;
		end
		32'h00001B94: begin
				q			<=			16'h00EF;
		end
		32'h00001B96: begin
				q			<=			16'h3C90;
		end
		32'h00001B98: begin
				q			<=			16'hA023;
		end
		32'h00001B9A: begin
				q			<=			16'hE2A9;
		end
		32'h00001B9C: begin
				q			<=			16'h1463;
		end
		32'h00001B9E: begin
				q			<=			16'h0405;
		end
		32'h00001BA0: begin
				q			<=			16'h0793;
		end
		32'h00001BA2: begin
				q			<=			16'hE244;
		end
		32'h00001BA4: begin
				q			<=			16'hC783;
		end
		32'h00001BA6: begin
				q			<=			16'h0097;
		end
		32'h00001BA8: begin
				q			<=			16'h8E63;
		end
		32'h00001BAA: begin
				q			<=			16'h0207;
		end
		32'h00001BAC: begin
				q			<=			16'h0793;
		end
		32'h00001BAE: begin
				q			<=			16'hE244;
		end
		32'h00001BB0: begin
				q			<=			16'hC783;
		end
		32'h00001BB2: begin
				q			<=			16'h0087;
		end
		32'h00001BB4: begin
				q			<=			16'hF793;
		end
		32'h00001BB6: begin
				q			<=			16'h0107;
		end
		32'h00001BB8: begin
				q			<=			16'h84E3;
		end
		32'h00001BBA: begin
				q			<=			16'hFA07;
		end
		32'h00001BBC: begin
				q			<=			16'h0693;
		end
		32'h00001BBE: begin
				q			<=			16'hE2DA;
		end
		32'h00001BC0: begin
				q			<=			16'h8613;
		end
		32'h00001BC2: begin
				q			<=			16'hD5CA;
		end
		32'h00001BC4: begin
				q			<=			16'h0593;
		end
		32'h00001BC6: begin
				q			<=			16'h1000;
		end
		32'h00001BC8: begin
				q			<=			16'h0513;
		end
		32'h00001BCA: begin
				q			<=			16'hD1C9;
		end
		32'h00001BCC: begin
				q			<=			16'h1097;
		end
		32'h00001BCE: begin
				q			<=			16'h0000;
		end
		32'h00001BD0: begin
				q			<=			16'h80E7;
		end
		32'h00001BD2: begin
				q			<=			16'h1A00;
		end
		32'h00001BD4: begin
				q			<=			16'h0593;
		end
		32'h00001BD6: begin
				q			<=			16'h0010;
		end
		32'h00001BD8: begin
				q			<=			16'h0513;
		end
		32'h00001BDA: begin
				q			<=			16'hD1C9;
		end
		32'h00001BDC: begin
				q			<=			16'hE0EF;
		end
		32'h00001BDE: begin
				q			<=			16'hFBDF;
		end
		32'h00001BE0: begin
				q			<=			16'hF06F;
		end
		32'h00001BE2: begin
				q			<=			16'hFA5F;
		end
		32'h00001BE4: begin
				q			<=			16'h2083;
		end
		32'h00001BE6: begin
				q			<=			16'h03C1;
		end
		32'h00001BE8: begin
				q			<=			16'h2403;
		end
		32'h00001BEA: begin
				q			<=			16'h0381;
		end
		32'h00001BEC: begin
				q			<=			16'h2483;
		end
		32'h00001BEE: begin
				q			<=			16'h0341;
		end
		32'h00001BF0: begin
				q			<=			16'h2903;
		end
		32'h00001BF2: begin
				q			<=			16'h0301;
		end
		32'h00001BF4: begin
				q			<=			16'h2983;
		end
		32'h00001BF6: begin
				q			<=			16'h02C1;
		end
		32'h00001BF8: begin
				q			<=			16'h2A03;
		end
		32'h00001BFA: begin
				q			<=			16'h0281;
		end
		32'h00001BFC: begin
				q			<=			16'h2A83;
		end
		32'h00001BFE: begin
				q			<=			16'h0241;
		end
		32'h00001C00: begin
				q			<=			16'h2B03;
		end
		32'h00001C02: begin
				q			<=			16'h0201;
		end
		32'h00001C04: begin
				q			<=			16'h0113;
		end
		32'h00001C06: begin
				q			<=			16'h0401;
		end
		32'h00001C08: begin
				q			<=			16'h8067;
		end
		32'h00001C0A: begin
				q			<=			16'h0000;
		end
		32'h00001C0C: begin
				q			<=			16'h0000;
		end
		32'h00001C0E: begin
				q			<=			16'h0000;
		end
		32'h00001C10: begin
				q			<=			16'h8067;
		end
		32'h00001C12: begin
				q			<=			16'h0000;
		end
		32'h00001C14: begin
				q			<=			16'h0000;
		end
		32'h00001C16: begin
				q			<=			16'h0000;
		end
		32'h00001C18: begin
				q			<=			16'h0513;
		end
		32'h00001C1A: begin
				q			<=			16'h0000;
		end
		32'h00001C1C: begin
				q			<=			16'h8067;
		end
		32'h00001C1E: begin
				q			<=			16'h0000;
		end
		32'h00001C20: begin
				q			<=			16'h0000;
		end
		32'h00001C22: begin
				q			<=			16'h0000;
		end
		32'h00001C24: begin
				q			<=			16'h0113;
		end
		32'h00001C26: begin
				q			<=			16'hFF01;
		end
		32'h00001C28: begin
				q			<=			16'h2623;
		end
		32'h00001C2A: begin
				q			<=			16'h0011;
		end
		32'h00001C2C: begin
				q			<=			16'h0313;
		end
		32'h00001C2E: begin
				q			<=			16'h0006;
		end
		32'h00001C30: begin
				q			<=			16'h17B7;
		end
		32'h00001C32: begin
				q			<=			16'h0001;
		end
		32'h00001C34: begin
				q			<=			16'hA783;
		end
		32'h00001C36: begin
				q			<=			16'h8F07;
		end
		32'h00001C38: begin
				q			<=			16'h8E63;
		end
		32'h00001C3A: begin
				q			<=			16'h04B7;
		end
		32'h00001C3C: begin
				q			<=			16'h07B7;
		end
		32'h00001C3E: begin
				q			<=			16'h8000;
		end
		32'h00001C40: begin
				q			<=			16'hA223;
		end
		32'h00001C42: begin
				q			<=			16'h00B7;
		end
		32'h00001C44: begin
				q			<=			16'h0713;
		end
		32'h00001C46: begin
				q			<=			16'h0010;
		end
		32'h00001C48: begin
				q			<=			16'hA423;
		end
		32'h00001C4A: begin
				q			<=			16'h00E7;
		end
		32'h00001C4C: begin
				q			<=			16'hA783;
		end
		32'h00001C4E: begin
				q			<=			16'h0087;
		end
		32'h00001C50: begin
				q			<=			16'hF793;
		end
		32'h00001C52: begin
				q			<=			16'h0087;
		end
		32'h00001C54: begin
				q			<=			16'h9263;
		end
		32'h00001C56: begin
				q			<=			16'h0607;
		end
		32'h00001C58: begin
				q			<=			16'h0737;
		end
		32'h00001C5A: begin
				q			<=			16'h8000;
		end
		32'h00001C5C: begin
				q			<=			16'h2783;
		end
		32'h00001C5E: begin
				q			<=			16'h0087;
		end
		32'h00001C60: begin
				q			<=			16'hF793;
		end
		32'h00001C62: begin
				q			<=			16'h0087;
		end
		32'h00001C64: begin
				q			<=			16'h8CE3;
		end
		32'h00001C66: begin
				q			<=			16'hFE07;
		end
		32'h00001C68: begin
				q			<=			16'h17B7;
		end
		32'h00001C6A: begin
				q			<=			16'h0001;
		end
		32'h00001C6C: begin
				q			<=			16'h8793;
		end
		32'h00001C6E: begin
				q			<=			16'h8F47;
		end
		32'h00001C70: begin
				q			<=			16'h08B7;
		end
		32'h00001C72: begin
				q			<=			16'h8000;
		end
		32'h00001C74: begin
				q			<=			16'h1837;
		end
		32'h00001C76: begin
				q			<=			16'h0001;
		end
		32'h00001C78: begin
				q			<=			16'h0813;
		end
		32'h00001C7A: begin
				q			<=			16'hAF48;
		end
		32'h00001C7C: begin
				q			<=			16'h8793;
		end
		32'h00001C7E: begin
				q			<=			16'h0047;
		end
		32'h00001C80: begin
				q			<=			16'hA703;
		end
		32'h00001C82: begin
				q			<=			16'h00C8;
		end
		32'h00001C84: begin
				q			<=			16'hAE23;
		end
		32'h00001C86: begin
				q			<=			16'hFEE7;
		end
		32'h00001C88: begin
				q			<=			16'h9AE3;
		end
		32'h00001C8A: begin
				q			<=			16'hFF07;
		end
		32'h00001C8C: begin
				q			<=			16'h17B7;
		end
		32'h00001C8E: begin
				q			<=			16'h0001;
		end
		32'h00001C90: begin
				q			<=			16'hA823;
		end
		32'h00001C92: begin
				q			<=			16'h8EB7;
		end
		32'h00001C94: begin
				q			<=			16'h8613;
		end
		32'h00001C96: begin
				q			<=			16'h0006;
		end
		32'h00001C98: begin
				q			<=			16'h17B7;
		end
		32'h00001C9A: begin
				q			<=			16'h0001;
		end
		32'h00001C9C: begin
				q			<=			16'h8793;
		end
		32'h00001C9E: begin
				q			<=			16'h8F47;
		end
		32'h00001CA0: begin
				q			<=			16'h85B3;
		end
		32'h00001CA2: begin
				q			<=			16'h0067;
		end
		32'h00001CA4: begin
				q			<=			16'h00EF;
		end
		32'h00001CA6: begin
				q			<=			16'h6550;
		end
		32'h00001CA8: begin
				q			<=			16'h0513;
		end
		32'h00001CAA: begin
				q			<=			16'h0000;
		end
		32'h00001CAC: begin
				q			<=			16'h2083;
		end
		32'h00001CAE: begin
				q			<=			16'h00C1;
		end
		32'h00001CB0: begin
				q			<=			16'h0113;
		end
		32'h00001CB2: begin
				q			<=			16'h0101;
		end
		32'h00001CB4: begin
				q			<=			16'h8067;
		end
		32'h00001CB6: begin
				q			<=			16'h0000;
		end
		32'h00001CB8: begin
				q			<=			16'h17B7;
		end
		32'h00001CBA: begin
				q			<=			16'h0001;
		end
		32'h00001CBC: begin
				q			<=			16'h8793;
		end
		32'h00001CBE: begin
				q			<=			16'h8F47;
		end
		32'h00001CC0: begin
				q			<=			16'hF06F;
		end
		32'h00001CC2: begin
				q			<=			16'hFB1F;
		end
		32'h00001CC4: begin
				q			<=			16'h0000;
		end
		32'h00001CC6: begin
				q			<=			16'h0000;
		end
		32'h00001CC8: begin
				q			<=			16'h4703;
		end
		32'h00001CCA: begin
				q			<=			16'h0035;
		end
		32'h00001CCC: begin
				q			<=			16'h1713;
		end
		32'h00001CCE: begin
				q			<=			16'h0087;
		end
		32'h00001CD0: begin
				q			<=			16'h4783;
		end
		32'h00001CD2: begin
				q			<=			16'h0025;
		end
		32'h00001CD4: begin
				q			<=			16'hE7B3;
		end
		32'h00001CD6: begin
				q			<=			16'h00E7;
		end
		32'h00001CD8: begin
				q			<=			16'h9713;
		end
		32'h00001CDA: begin
				q			<=			16'h0087;
		end
		32'h00001CDC: begin
				q			<=			16'h4783;
		end
		32'h00001CDE: begin
				q			<=			16'h0015;
		end
		32'h00001CE0: begin
				q			<=			16'hE7B3;
		end
		32'h00001CE2: begin
				q			<=			16'h00E7;
		end
		32'h00001CE4: begin
				q			<=			16'h9793;
		end
		32'h00001CE6: begin
				q			<=			16'h0087;
		end
		32'h00001CE8: begin
				q			<=			16'h4503;
		end
		32'h00001CEA: begin
				q			<=			16'h0005;
		end
		32'h00001CEC: begin
				q			<=			16'h6533;
		end
		32'h00001CEE: begin
				q			<=			16'h00F5;
		end
		32'h00001CF0: begin
				q			<=			16'h8067;
		end
		32'h00001CF2: begin
				q			<=			16'h0000;
		end
		32'h00001CF4: begin
				q			<=			16'h0000;
		end
		32'h00001CF6: begin
				q			<=			16'h0000;
		end
		32'h00001CF8: begin
				q			<=			16'h17B7;
		end
		32'h00001CFA: begin
				q			<=			16'h0001;
		end
		32'h00001CFC: begin
				q			<=			16'hA703;
		end
		32'h00001CFE: begin
				q			<=			16'hF9C7;
		end
		32'h00001D00: begin
				q			<=			16'h0693;
		end
		32'h00001D02: begin
				q			<=			16'hFFE5;
		end
		32'h00001D04: begin
				q			<=			16'h2783;
		end
		32'h00001D06: begin
				q			<=			16'h0087;
		end
		32'h00001D08: begin
				q			<=			16'h8793;
		end
		32'h00001D0A: begin
				q			<=			16'hFFE7;
		end
		32'h00001D0C: begin
				q			<=			16'hFC63;
		end
		32'h00001D0E: begin
				q			<=			16'h00F6;
		end
		32'h00001D10: begin
				q			<=			16'h4503;
		end
		32'h00001D12: begin
				q			<=			16'h0027;
		end
		32'h00001D14: begin
				q			<=			16'h0533;
		end
		32'h00001D16: begin
				q			<=			16'h02D5;
		end
		32'h00001D18: begin
				q			<=			16'h2783;
		end
		32'h00001D1A: begin
				q			<=			16'h0147;
		end
		32'h00001D1C: begin
				q			<=			16'h0533;
		end
		32'h00001D1E: begin
				q			<=			16'h00F5;
		end
		32'h00001D20: begin
				q			<=			16'h8067;
		end
		32'h00001D22: begin
				q			<=			16'h0000;
		end
		32'h00001D24: begin
				q			<=			16'h0513;
		end
		32'h00001D26: begin
				q			<=			16'h0000;
		end
		32'h00001D28: begin
				q			<=			16'h8067;
		end
		32'h00001D2A: begin
				q			<=			16'h0000;
		end
		32'h00001D2C: begin
				q			<=			16'h0000;
		end
		32'h00001D2E: begin
				q			<=			16'h0000;
		end
		32'h00001D30: begin
				q			<=			16'h1737;
		end
		32'h00001D32: begin
				q			<=			16'h0001;
		end
		32'h00001D34: begin
				q			<=			16'h2683;
		end
		32'h00001D36: begin
				q			<=			16'hF9C7;
		end
		32'h00001D38: begin
				q			<=			16'h1023;
		end
		32'h00001D3A: begin
				q			<=			16'h0005;
		end
		32'h00001D3C: begin
				q			<=			16'h2703;
		end
		32'h00001D3E: begin
				q			<=			16'h0085;
		end
		32'h00001D40: begin
				q			<=			16'h0613;
		end
		32'h00001D42: begin
				q			<=			16'h0010;
		end
		32'h00001D44: begin
				q			<=			16'h0663;
		end
		32'h00001D46: begin
				q			<=			16'h04C7;
		end
		32'h00001D48: begin
				q			<=			16'h0113;
		end
		32'h00001D4A: begin
				q			<=			16'hFF01;
		end
		32'h00001D4C: begin
				q			<=			16'h2623;
		end
		32'h00001D4E: begin
				q			<=			16'h0011;
		end
		32'h00001D50: begin
				q			<=			16'h2423;
		end
		32'h00001D52: begin
				q			<=			16'h0081;
		end
		32'h00001D54: begin
				q			<=			16'h0413;
		end
		32'h00001D56: begin
				q			<=			16'h0005;
		end
		32'h00001D58: begin
				q			<=			16'hA603;
		end
		32'h00001D5A: begin
				q			<=			16'h0086;
		end
		32'h00001D5C: begin
				q			<=			16'h0513;
		end
		32'h00001D5E: begin
				q			<=			16'h0010;
		end
		32'h00001D60: begin
				q			<=			16'h7663;
		end
		32'h00001D62: begin
				q			<=			16'h04C7;
		end
		32'h00001D64: begin
				q			<=			16'h1A63;
		end
		32'h00001D66: begin
				q			<=			16'h0207;
		end
		32'h00001D68: begin
				q			<=			16'hC703;
		end
		32'h00001D6A: begin
				q			<=			16'h0006;
		end
		32'h00001D6C: begin
				q			<=			16'h0793;
		end
		32'h00001D6E: begin
				q			<=			16'h0030;
		end
		32'h00001D70: begin
				q			<=			16'h0863;
		end
		32'h00001D72: begin
				q			<=			16'h00F7;
		end
		32'h00001D74: begin
				q			<=			16'h2623;
		end
		32'h00001D76: begin
				q			<=			16'h0004;
		end
		32'h00001D78: begin
				q			<=			16'hA503;
		end
		32'h00001D7A: begin
				q			<=			16'h0106;
		end
		32'h00001D7C: begin
				q			<=			16'h006F;
		end
		32'h00001D7E: begin
				q			<=			16'h0280;
		end
		32'h00001D80: begin
				q			<=			16'hA703;
		end
		32'h00001D82: begin
				q			<=			16'h0106;
		end
		32'h00001D84: begin
				q			<=			16'h2623;
		end
		32'h00001D86: begin
				q			<=			16'h00E4;
		end
		32'h00001D88: begin
				q			<=			16'h08E3;
		end
		32'h00001D8A: begin
				q			<=			16'hFE07;
		end
		32'h00001D8C: begin
				q			<=			16'h006F;
		end
		32'h00001D8E: begin
				q			<=			16'h0100;
		end
		32'h00001D90: begin
				q			<=			16'h0513;
		end
		32'h00001D92: begin
				q			<=			16'h0010;
		end
		32'h00001D94: begin
				q			<=			16'h8067;
		end
		32'h00001D96: begin
				q			<=			16'h0000;
		end
		32'h00001D98: begin
				q			<=			16'h2623;
		end
		32'h00001D9A: begin
				q			<=			16'h00E4;
		end
		32'h00001D9C: begin
				q			<=			16'h0513;
		end
		32'h00001D9E: begin
				q			<=			16'h0007;
		end
		32'h00001DA0: begin
				q			<=			16'hF0EF;
		end
		32'h00001DA2: begin
				q			<=			16'hF59F;
		end
		32'h00001DA4: begin
				q			<=			16'h2823;
		end
		32'h00001DA6: begin
				q			<=			16'h00A4;
		end
		32'h00001DA8: begin
				q			<=			16'h0513;
		end
		32'h00001DAA: begin
				q			<=			16'h0000;
		end
		32'h00001DAC: begin
				q			<=			16'h2083;
		end
		32'h00001DAE: begin
				q			<=			16'h00C1;
		end
		32'h00001DB0: begin
				q			<=			16'h2403;
		end
		32'h00001DB2: begin
				q			<=			16'h0081;
		end
		32'h00001DB4: begin
				q			<=			16'h0113;
		end
		32'h00001DB6: begin
				q			<=			16'h0101;
		end
		32'h00001DB8: begin
				q			<=			16'h8067;
		end
		32'h00001DBA: begin
				q			<=			16'h0000;
		end
		32'h00001DBC: begin
				q			<=			16'h0000;
		end
		32'h00001DBE: begin
				q			<=			16'h0000;
		end
		32'h00001DC0: begin
				q			<=			16'h0793;
		end
		32'h00001DC2: begin
				q			<=			16'h0010;
		end
		32'h00001DC4: begin
				q			<=			16'hF263;
		end
		32'h00001DC6: begin
				q			<=			16'h0CA7;
		end
		32'h00001DC8: begin
				q			<=			16'h17B7;
		end
		32'h00001DCA: begin
				q			<=			16'h0001;
		end
		32'h00001DCC: begin
				q			<=			16'hA703;
		end
		32'h00001DCE: begin
				q			<=			16'hF9C7;
		end
		32'h00001DD0: begin
				q			<=			16'h2683;
		end
		32'h00001DD2: begin
				q			<=			16'h0087;
		end
		32'h00001DD4: begin
				q			<=			16'h0793;
		end
		32'h00001DD6: begin
				q			<=			16'h0010;
		end
		32'h00001DD8: begin
				q			<=			16'h7A63;
		end
		32'h00001DDA: begin
				q			<=			16'h0AD5;
		end
		32'h00001DDC: begin
				q			<=			16'h0113;
		end
		32'h00001DDE: begin
				q			<=			16'hFE01;
		end
		32'h00001DE0: begin
				q			<=			16'h2E23;
		end
		32'h00001DE2: begin
				q			<=			16'h0011;
		end
		32'h00001DE4: begin
				q			<=			16'h4783;
		end
		32'h00001DE6: begin
				q			<=			16'h0007;
		end
		32'h00001DE8: begin
				q			<=			16'h0693;
		end
		32'h00001DEA: begin
				q			<=			16'h0020;
		end
		32'h00001DEC: begin
				q			<=			16'h8063;
		end
		32'h00001DEE: begin
				q			<=			16'h02D7;
		end
		32'h00001DF0: begin
				q			<=			16'h0693;
		end
		32'h00001DF2: begin
				q			<=			16'h0030;
		end
		32'h00001DF4: begin
				q			<=			16'h8A63;
		end
		32'h00001DF6: begin
				q			<=			16'h04D7;
		end
		32'h00001DF8: begin
				q			<=			16'h0793;
		end
		32'h00001DFA: begin
				q			<=			16'h0010;
		end
		32'h00001DFC: begin
				q			<=			16'h8513;
		end
		32'h00001DFE: begin
				q			<=			16'h0007;
		end
		32'h00001E00: begin
				q			<=			16'h2083;
		end
		32'h00001E02: begin
				q			<=			16'h01C1;
		end
		32'h00001E04: begin
				q			<=			16'h0113;
		end
		32'h00001E06: begin
				q			<=			16'h0201;
		end
		32'h00001E08: begin
				q			<=			16'h8067;
		end
		32'h00001E0A: begin
				q			<=			16'h0000;
		end
		32'h00001E0C: begin
				q			<=			16'h7613;
		end
		32'h00001E0E: begin
				q			<=			16'h0FF5;
		end
		32'h00001E10: begin
				q			<=			16'h5513;
		end
		32'h00001E12: begin
				q			<=			16'h0085;
		end
		32'h00001E14: begin
				q			<=			16'h2583;
		end
		32'h00001E16: begin
				q			<=			16'h00C7;
		end
		32'h00001E18: begin
				q			<=			16'h0693;
		end
		32'h00001E1A: begin
				q			<=			16'h0020;
		end
		32'h00001E1C: begin
				q			<=			16'h1613;
		end
		32'h00001E1E: begin
				q			<=			16'h0016;
		end
		32'h00001E20: begin
				q			<=			16'h05B3;
		end
		32'h00001E22: begin
				q			<=			16'h00B5;
		end
		32'h00001E24: begin
				q			<=			16'h0513;
		end
		32'h00001E26: begin
				q			<=			16'h00C1;
		end
		32'h00001E28: begin
				q			<=			16'hF0EF;
		end
		32'h00001E2A: begin
				q			<=			16'hDFDF;
		end
		32'h00001E2C: begin
				q			<=			16'h0793;
		end
		32'h00001E2E: begin
				q			<=			16'h0010;
		end
		32'h00001E30: begin
				q			<=			16'h16E3;
		end
		32'h00001E32: begin
				q			<=			16'hFC05;
		end
		32'h00001E34: begin
				q			<=			16'h4783;
		end
		32'h00001E36: begin
				q			<=			16'h00D1;
		end
		32'h00001E38: begin
				q			<=			16'h9793;
		end
		32'h00001E3A: begin
				q			<=			16'h0087;
		end
		32'h00001E3C: begin
				q			<=			16'h4703;
		end
		32'h00001E3E: begin
				q			<=			16'h00C1;
		end
		32'h00001E40: begin
				q			<=			16'hE7B3;
		end
		32'h00001E42: begin
				q			<=			16'h00E7;
		end
		32'h00001E44: begin
				q			<=			16'hF06F;
		end
		32'h00001E46: begin
				q			<=			16'hFB9F;
		end
		32'h00001E48: begin
				q			<=			16'h7613;
		end
		32'h00001E4A: begin
				q			<=			16'h07F5;
		end
		32'h00001E4C: begin
				q			<=			16'h5513;
		end
		32'h00001E4E: begin
				q			<=			16'h0075;
		end
		32'h00001E50: begin
				q			<=			16'h2583;
		end
		32'h00001E52: begin
				q			<=			16'h00C7;
		end
		32'h00001E54: begin
				q			<=			16'h0693;
		end
		32'h00001E56: begin
				q			<=			16'h0040;
		end
		32'h00001E58: begin
				q			<=			16'h1613;
		end
		32'h00001E5A: begin
				q			<=			16'h0026;
		end
		32'h00001E5C: begin
				q			<=			16'h05B3;
		end
		32'h00001E5E: begin
				q			<=			16'h00B5;
		end
		32'h00001E60: begin
				q			<=			16'h0513;
		end
		32'h00001E62: begin
				q			<=			16'h00C1;
		end
		32'h00001E64: begin
				q			<=			16'hF0EF;
		end
		32'h00001E66: begin
				q			<=			16'hDC1F;
		end
		32'h00001E68: begin
				q			<=			16'h0793;
		end
		32'h00001E6A: begin
				q			<=			16'h0010;
		end
		32'h00001E6C: begin
				q			<=			16'h18E3;
		end
		32'h00001E6E: begin
				q			<=			16'hF805;
		end
		32'h00001E70: begin
				q			<=			16'h0513;
		end
		32'h00001E72: begin
				q			<=			16'h00C1;
		end
		32'h00001E74: begin
				q			<=			16'hF0EF;
		end
		32'h00001E76: begin
				q			<=			16'hE55F;
		end
		32'h00001E78: begin
				q			<=			16'h07B7;
		end
		32'h00001E7A: begin
				q			<=			16'h1000;
		end
		32'h00001E7C: begin
				q			<=			16'h8793;
		end
		32'h00001E7E: begin
				q			<=			16'hFFF7;
		end
		32'h00001E80: begin
				q			<=			16'h77B3;
		end
		32'h00001E82: begin
				q			<=			16'h00F5;
		end
		32'h00001E84: begin
				q			<=			16'hF06F;
		end
		32'h00001E86: begin
				q			<=			16'hF79F;
		end
		32'h00001E88: begin
				q			<=			16'h0793;
		end
		32'h00001E8A: begin
				q			<=			16'h0010;
		end
		32'h00001E8C: begin
				q			<=			16'h8513;
		end
		32'h00001E8E: begin
				q			<=			16'h0007;
		end
		32'h00001E90: begin
				q			<=			16'h8067;
		end
		32'h00001E92: begin
				q			<=			16'h0000;
		end
		32'h00001E94: begin
				q			<=			16'h0000;
		end
		32'h00001E96: begin
				q			<=			16'h0000;
		end
		32'h00001E98: begin
				q			<=			16'h0113;
		end
		32'h00001E9A: begin
				q			<=			16'hFF01;
		end
		32'h00001E9C: begin
				q			<=			16'h2623;
		end
		32'h00001E9E: begin
				q			<=			16'h0011;
		end
		32'h00001EA0: begin
				q			<=			16'h2423;
		end
		32'h00001EA2: begin
				q			<=			16'h0081;
		end
		32'h00001EA4: begin
				q			<=			16'h2223;
		end
		32'h00001EA6: begin
				q			<=			16'h0091;
		end
		32'h00001EA8: begin
				q			<=			16'h2023;
		end
		32'h00001EAA: begin
				q			<=			16'h0121;
		end
		32'h00001EAC: begin
				q			<=			16'h5403;
		end
		32'h00001EAE: begin
				q			<=			16'h0005;
		end
		32'h00001EB0: begin
				q			<=			16'h0413;
		end
		32'h00001EB2: begin
				q			<=			16'h0014;
		end
		32'h00001EB4: begin
				q			<=			16'h1413;
		end
		32'h00001EB6: begin
				q			<=			16'h0104;
		end
		32'h00001EB8: begin
				q			<=			16'h5413;
		end
		32'h00001EBA: begin
				q			<=			16'h0104;
		end
		32'h00001EBC: begin
				q			<=			16'h0793;
		end
		32'h00001EBE: begin
				q			<=			16'h0030;
		end
		32'h00001EC0: begin
				q			<=			16'h0463;
		end
		32'h00001EC2: begin
				q			<=			16'h0404;
		end
		32'h00001EC4: begin
				q			<=			16'h2703;
		end
		32'h00001EC6: begin
				q			<=			16'h0105;
		end
		32'h00001EC8: begin
				q			<=			16'h0793;
		end
		32'h00001ECA: begin
				q			<=			16'h0030;
		end
		32'h00001ECC: begin
				q			<=			16'h0E63;
		end
		32'h00001ECE: begin
				q			<=			16'h0207;
		end
		32'h00001ED0: begin
				q			<=			16'h0493;
		end
		32'h00001ED2: begin
				q			<=			16'h0005;
		end
		32'h00001ED4: begin
				q			<=			16'h7793;
		end
		32'h00001ED6: begin
				q			<=			16'h00F4;
		end
		32'h00001ED8: begin
				q			<=			16'h9463;
		end
		32'h00001EDA: begin
				q			<=			16'h0207;
		end
		32'h00001EDC: begin
				q			<=			16'h17B7;
		end
		32'h00001EDE: begin
				q			<=			16'h0001;
		end
		32'h00001EE0: begin
				q			<=			16'hA903;
		end
		32'h00001EE2: begin
				q			<=			16'hF9C7;
		end
		32'h00001EE4: begin
				q			<=			16'h0713;
		end
		32'h00001EE6: begin
				q			<=			16'h0017;
		end
		32'h00001EE8: begin
				q			<=			16'h2823;
		end
		32'h00001EEA: begin
				q			<=			16'h00E5;
		end
		32'h00001EEC: begin
				q			<=			16'h2503;
		end
		32'h00001EEE: begin
				q			<=			16'h00C5;
		end
		32'h00001EF0: begin
				q			<=			16'h1A63;
		end
		32'h00001EF2: begin
				q			<=			16'h0205;
		end
		32'h00001EF4: begin
				q			<=			16'h5703;
		end
		32'h00001EF6: begin
				q			<=			16'h0049;
		end
		32'h00001EF8: begin
				q			<=			16'h0793;
		end
		32'h00001EFA: begin
				q			<=			16'h0030;
		end
		32'h00001EFC: begin
				q			<=			16'h7663;
		end
		32'h00001EFE: begin
				q			<=			16'h00E4;
		end
		32'h00001F00: begin
				q			<=			16'h9023;
		end
		32'h00001F02: begin
				q			<=			16'h0084;
		end
		32'h00001F04: begin
				q			<=			16'h0793;
		end
		32'h00001F06: begin
				q			<=			16'h0000;
		end
		32'h00001F08: begin
				q			<=			16'h8513;
		end
		32'h00001F0A: begin
				q			<=			16'h0007;
		end
		32'h00001F0C: begin
				q			<=			16'h2083;
		end
		32'h00001F0E: begin
				q			<=			16'h00C1;
		end
		32'h00001F10: begin
				q			<=			16'h2403;
		end
		32'h00001F12: begin
				q			<=			16'h0081;
		end
		32'h00001F14: begin
				q			<=			16'h2483;
		end
		32'h00001F16: begin
				q			<=			16'h0041;
		end
		32'h00001F18: begin
				q			<=			16'h2903;
		end
		32'h00001F1A: begin
				q			<=			16'h0001;
		end
		32'h00001F1C: begin
				q			<=			16'h0113;
		end
		32'h00001F1E: begin
				q			<=			16'h0101;
		end
		32'h00001F20: begin
				q			<=			16'h8067;
		end
		32'h00001F22: begin
				q			<=			16'h0000;
		end
		32'h00001F24: begin
				q			<=			16'h4783;
		end
		32'h00001F26: begin
				q			<=			16'h0029;
		end
		32'h00001F28: begin
				q			<=			16'h8793;
		end
		32'h00001F2A: begin
				q			<=			16'hFFF7;
		end
		32'h00001F2C: begin
				q			<=			16'h5713;
		end
		32'h00001F2E: begin
				q			<=			16'h0044;
		end
		32'h00001F30: begin
				q			<=			16'hF7B3;
		end
		32'h00001F32: begin
				q			<=			16'h00E7;
		end
		32'h00001F34: begin
				q			<=			16'h96E3;
		end
		32'h00001F36: begin
				q			<=			16'hFC07;
		end
		32'h00001F38: begin
				q			<=			16'hF0EF;
		end
		32'h00001F3A: begin
				q			<=			16'hE89F;
		end
		32'h00001F3C: begin
				q			<=			16'h0713;
		end
		32'h00001F3E: begin
				q			<=			16'h0010;
		end
		32'h00001F40: begin
				q			<=			16'h0793;
		end
		32'h00001F42: begin
				q			<=			16'h0010;
		end
		32'h00001F44: begin
				q			<=			16'h72E3;
		end
		32'h00001F46: begin
				q			<=			16'hFCA7;
		end
		32'h00001F48: begin
				q			<=			16'h2703;
		end
		32'h00001F4A: begin
				q			<=			16'h0089;
		end
		32'h00001F4C: begin
				q			<=			16'h0793;
		end
		32'h00001F4E: begin
				q			<=			16'h0030;
		end
		32'h00001F50: begin
				q			<=			16'h7CE3;
		end
		32'h00001F52: begin
				q			<=			16'hFAE5;
		end
		32'h00001F54: begin
				q			<=			16'hA623;
		end
		32'h00001F56: begin
				q			<=			16'h00A4;
		end
		32'h00001F58: begin
				q			<=			16'hF0EF;
		end
		32'h00001F5A: begin
				q			<=			16'hDA1F;
		end
		32'h00001F5C: begin
				q			<=			16'hA823;
		end
		32'h00001F5E: begin
				q			<=			16'h00A4;
		end
		32'h00001F60: begin
				q			<=			16'hF06F;
		end
		32'h00001F62: begin
				q			<=			16'hFA1F;
		end
		32'h00001F64: begin
				q			<=			16'h0000;
		end
		32'h00001F66: begin
				q			<=			16'h0000;
		end
		32'h00001F68: begin
				q			<=			16'h0113;
		end
		32'h00001F6A: begin
				q			<=			16'hFF01;
		end
		32'h00001F6C: begin
				q			<=			16'h2623;
		end
		32'h00001F6E: begin
				q			<=			16'h0011;
		end
		32'h00001F70: begin
				q			<=			16'h2423;
		end
		32'h00001F72: begin
				q			<=			16'h0081;
		end
		32'h00001F74: begin
				q			<=			16'h2223;
		end
		32'h00001F76: begin
				q			<=			16'h0091;
		end
		32'h00001F78: begin
				q			<=			16'h0413;
		end
		32'h00001F7A: begin
				q			<=			16'h0005;
		end
		32'h00001F7C: begin
				q			<=			16'h8493;
		end
		32'h00001F7E: begin
				q			<=			16'h0005;
		end
		32'h00001F80: begin
				q			<=			16'h0693;
		end
		32'h00001F82: begin
				q			<=			16'h0020;
		end
		32'h00001F84: begin
				q			<=			16'h0613;
		end
		32'h00001F86: begin
				q			<=			16'h1FE0;
		end
		32'h00001F88: begin
				q			<=			16'hF0EF;
		end
		32'h00001F8A: begin
				q			<=			16'hC9DF;
		end
		32'h00001F8C: begin
				q			<=			16'h0713;
		end
		32'h00001F8E: begin
				q			<=			16'h0030;
		end
		32'h00001F90: begin
				q			<=			16'h1663;
		end
		32'h00001F92: begin
				q			<=			16'h0205;
		end
		32'h00001F94: begin
				q			<=			16'h4783;
		end
		32'h00001F96: begin
				q			<=			16'h0014;
		end
		32'h00001F98: begin
				q			<=			16'h9793;
		end
		32'h00001F9A: begin
				q			<=			16'h0087;
		end
		32'h00001F9C: begin
				q			<=			16'h4703;
		end
		32'h00001F9E: begin
				q			<=			16'h0004;
		end
		32'h00001FA0: begin
				q			<=			16'hE7B3;
		end
		32'h00001FA2: begin
				q			<=			16'h00E7;
		end
		32'h00001FA4: begin
				q			<=			16'h9793;
		end
		32'h00001FA6: begin
				q			<=			16'h0107;
		end
		32'h00001FA8: begin
				q			<=			16'hD793;
		end
		32'h00001FAA: begin
				q			<=			16'h4107;
		end
		32'h00001FAC: begin
				q			<=			16'hB6B7;
		end
		32'h00001FAE: begin
				q			<=			16'hFFFF;
		end
		32'h00001FB0: begin
				q			<=			16'h8693;
		end
		32'h00001FB2: begin
				q			<=			16'hA556;
		end
		32'h00001FB4: begin
				q			<=			16'h0713;
		end
		32'h00001FB6: begin
				q			<=			16'h0020;
		end
		32'h00001FB8: begin
				q			<=			16'h8E63;
		end
		32'h00001FBA: begin
				q			<=			16'h00D7;
		end
		32'h00001FBC: begin
				q			<=			16'h0513;
		end
		32'h00001FBE: begin
				q			<=			16'h0007;
		end
		32'h00001FC0: begin
				q			<=			16'h2083;
		end
		32'h00001FC2: begin
				q			<=			16'h00C1;
		end
		32'h00001FC4: begin
				q			<=			16'h2403;
		end
		32'h00001FC6: begin
				q			<=			16'h0081;
		end
		32'h00001FC8: begin
				q			<=			16'h2483;
		end
		32'h00001FCA: begin
				q			<=			16'h0041;
		end
		32'h00001FCC: begin
				q			<=			16'h0113;
		end
		32'h00001FCE: begin
				q			<=			16'h0101;
		end
		32'h00001FD0: begin
				q			<=			16'h8067;
		end
		32'h00001FD2: begin
				q			<=			16'h0000;
		end
		32'h00001FD4: begin
				q			<=			16'h0693;
		end
		32'h00001FD6: begin
				q			<=			16'h0020;
		end
		32'h00001FD8: begin
				q			<=			16'h0613;
		end
		32'h00001FDA: begin
				q			<=			16'h0360;
		end
		32'h00001FDC: begin
				q			<=			16'h8593;
		end
		32'h00001FDE: begin
				q			<=			16'h0004;
		end
		32'h00001FE0: begin
				q			<=			16'h0513;
		end
		32'h00001FE2: begin
				q			<=			16'h0004;
		end
		32'h00001FE4: begin
				q			<=			16'hF0EF;
		end
		32'h00001FE6: begin
				q			<=			16'hC41F;
		end
		32'h00001FE8: begin
				q			<=			16'h1663;
		end
		32'h00001FEA: begin
				q			<=			16'h0205;
		end
		32'h00001FEC: begin
				q			<=			16'h4783;
		end
		32'h00001FEE: begin
				q			<=			16'h0014;
		end
		32'h00001FF0: begin
				q			<=			16'h9793;
		end
		32'h00001FF2: begin
				q			<=			16'h0087;
		end
		32'h00001FF4: begin
				q			<=			16'h4703;
		end
		32'h00001FF6: begin
				q			<=			16'h0004;
		end
		32'h00001FF8: begin
				q			<=			16'hE7B3;
		end
		32'h00001FFA: begin
				q			<=			16'h00E7;
		end
		32'h00001FFC: begin
				q			<=			16'h9793;
		end
		32'h00001FFE: begin
				q			<=			16'h0107;
		end
		32'h00002000: begin
				q			<=			16'hD793;
		end
		32'h00002002: begin
				q			<=			16'h4107;
		end
		32'h00002004: begin
				q			<=			16'h46B7;
		end
		32'h00002006: begin
				q			<=			16'h0000;
		end
		32'h00002008: begin
				q			<=			16'h8693;
		end
		32'h0000200A: begin
				q			<=			16'h1466;
		end
		32'h0000200C: begin
				q			<=			16'h0713;
		end
		32'h0000200E: begin
				q			<=			16'h0000;
		end
		32'h00002010: begin
				q			<=			16'h86E3;
		end
		32'h00002012: begin
				q			<=			16'hFAD7;
		end
		32'h00002014: begin
				q			<=			16'h0693;
		end
		32'h00002016: begin
				q			<=			16'h0020;
		end
		32'h00002018: begin
				q			<=			16'h0613;
		end
		32'h0000201A: begin
				q			<=			16'h0520;
		end
		32'h0000201C: begin
				q			<=			16'h8593;
		end
		32'h0000201E: begin
				q			<=			16'h0004;
		end
		32'h00002020: begin
				q			<=			16'h0513;
		end
		32'h00002022: begin
				q			<=			16'h0004;
		end
		32'h00002024: begin
				q			<=			16'hF0EF;
		end
		32'h00002026: begin
				q			<=			16'hC01F;
		end
		32'h00002028: begin
				q			<=			16'h0713;
		end
		32'h0000202A: begin
				q			<=			16'h0010;
		end
		32'h0000202C: begin
				q			<=			16'h18E3;
		end
		32'h0000202E: begin
				q			<=			16'hF805;
		end
		32'h00002030: begin
				q			<=			16'h4703;
		end
		32'h00002032: begin
				q			<=			16'h0014;
		end
		32'h00002034: begin
				q			<=			16'h1713;
		end
		32'h00002036: begin
				q			<=			16'h0087;
		end
		32'h00002038: begin
				q			<=			16'h4783;
		end
		32'h0000203A: begin
				q			<=			16'h0004;
		end
		32'h0000203C: begin
				q			<=			16'h6733;
		end
		32'h0000203E: begin
				q			<=			16'h00F7;
		end
		32'h00002040: begin
				q			<=			16'h1713;
		end
		32'h00002042: begin
				q			<=			16'h0107;
		end
		32'h00002044: begin
				q			<=			16'h5713;
		end
		32'h00002046: begin
				q			<=			16'h4107;
		end
		32'h00002048: begin
				q			<=			16'hC7B7;
		end
		32'h0000204A: begin
				q			<=			16'hFFFF;
		end
		32'h0000204C: begin
				q			<=			16'h8793;
		end
		32'h0000204E: begin
				q			<=			16'hEBA7;
		end
		32'h00002050: begin
				q			<=			16'h0733;
		end
		32'h00002052: begin
				q			<=			16'h00F7;
		end
		32'h00002054: begin
				q			<=			16'h3733;
		end
		32'h00002056: begin
				q			<=			16'h00E0;
		end
		32'h00002058: begin
				q			<=			16'hF06F;
		end
		32'h0000205A: begin
				q			<=			16'hF65F;
		end
		32'h0000205C: begin
				q			<=			16'h0000;
		end
		32'h0000205E: begin
				q			<=			16'h0000;
		end
		32'h00002060: begin
				q			<=			16'h17B7;
		end
		32'h00002062: begin
				q			<=			16'h0001;
		end
		32'h00002064: begin
				q			<=			16'hA783;
		end
		32'h00002066: begin
				q			<=			16'hF9C7;
		end
		32'h00002068: begin
				q			<=			16'hC703;
		end
		32'h0000206A: begin
				q			<=			16'h0007;
		end
		32'h0000206C: begin
				q			<=			16'h0793;
		end
		32'h0000206E: begin
				q			<=			16'h0030;
		end
		32'h00002070: begin
				q			<=			16'h0063;
		end
		32'h00002072: begin
				q			<=			16'h02F7;
		end
		32'h00002074: begin
				q			<=			16'h0713;
		end
		32'h00002076: begin
				q			<=			16'h0000;
		end
		32'h00002078: begin
				q			<=			16'h4783;
		end
		32'h0000207A: begin
				q			<=			16'h01B5;
		end
		32'h0000207C: begin
				q			<=			16'h9793;
		end
		32'h0000207E: begin
				q			<=			16'h0087;
		end
		32'h00002080: begin
				q			<=			16'h4503;
		end
		32'h00002082: begin
				q			<=			16'h01A5;
		end
		32'h00002084: begin
				q			<=			16'hE533;
		end
		32'h00002086: begin
				q			<=			16'h00A7;
		end
		32'h00002088: begin
				q			<=			16'h6533;
		end
		32'h0000208A: begin
				q			<=			16'h00E5;
		end
		32'h0000208C: begin
				q			<=			16'h8067;
		end
		32'h0000208E: begin
				q			<=			16'h0000;
		end
		32'h00002090: begin
				q			<=			16'h4703;
		end
		32'h00002092: begin
				q			<=			16'h0155;
		end
		32'h00002094: begin
				q			<=			16'h1713;
		end
		32'h00002096: begin
				q			<=			16'h0087;
		end
		32'h00002098: begin
				q			<=			16'h4783;
		end
		32'h0000209A: begin
				q			<=			16'h0145;
		end
		32'h0000209C: begin
				q			<=			16'h6733;
		end
		32'h0000209E: begin
				q			<=			16'h00F7;
		end
		32'h000020A0: begin
				q			<=			16'h1713;
		end
		32'h000020A2: begin
				q			<=			16'h0107;
		end
		32'h000020A4: begin
				q			<=			16'hF06F;
		end
		32'h000020A6: begin
				q			<=			16'hFD5F;
		end
		32'h000020A8: begin
				q			<=			16'h0000;
		end
		32'h000020AA: begin
				q			<=			16'h0000;
		end
		32'h000020AC: begin
				q			<=			16'h0113;
		end
		32'h000020AE: begin
				q			<=			16'hFD01;
		end
		32'h000020B0: begin
				q			<=			16'h2623;
		end
		32'h000020B2: begin
				q			<=			16'h0211;
		end
		32'h000020B4: begin
				q			<=			16'h2423;
		end
		32'h000020B6: begin
				q			<=			16'h0281;
		end
		32'h000020B8: begin
				q			<=			16'h2223;
		end
		32'h000020BA: begin
				q			<=			16'h0291;
		end
		32'h000020BC: begin
				q			<=			16'h2023;
		end
		32'h000020BE: begin
				q			<=			16'h0321;
		end
		32'h000020C0: begin
				q			<=			16'h2E23;
		end
		32'h000020C2: begin
				q			<=			16'h0131;
		end
		32'h000020C4: begin
				q			<=			16'h2C23;
		end
		32'h000020C6: begin
				q			<=			16'h0141;
		end
		32'h000020C8: begin
				q			<=			16'h2A23;
		end
		32'h000020CA: begin
				q			<=			16'h0151;
		end
		32'h000020CC: begin
				q			<=			16'h2823;
		end
		32'h000020CE: begin
				q			<=			16'h0161;
		end
		32'h000020D0: begin
				q			<=			16'h2623;
		end
		32'h000020D2: begin
				q			<=			16'h0171;
		end
		32'h000020D4: begin
				q			<=			16'h2423;
		end
		32'h000020D6: begin
				q			<=			16'h0181;
		end
		32'h000020D8: begin
				q			<=			16'h0413;
		end
		32'h000020DA: begin
				q			<=			16'h0005;
		end
		32'h000020DC: begin
				q			<=			16'h8493;
		end
		32'h000020DE: begin
				q			<=			16'h0005;
		end
		32'h000020E0: begin
				q			<=			16'h0913;
		end
		32'h000020E2: begin
				q			<=			16'h0006;
		end
		32'h000020E4: begin
				q			<=			16'h4783;
		end
		32'h000020E6: begin
				q			<=			16'h0006;
		end
		32'h000020E8: begin
				q			<=			16'h0713;
		end
		32'h000020EA: begin
				q			<=			16'h0200;
		end
		32'h000020EC: begin
				q			<=			16'h9863;
		end
		32'h000020EE: begin
				q			<=			16'h00E7;
		end
		32'h000020F0: begin
				q			<=			16'h0913;
		end
		32'h000020F2: begin
				q			<=			16'h0019;
		end
		32'h000020F4: begin
				q			<=			16'h4783;
		end
		32'h000020F6: begin
				q			<=			16'h0009;
		end
		32'h000020F8: begin
				q			<=			16'h8CE3;
		end
		32'h000020FA: begin
				q			<=			16'hFEE7;
		end
		32'h000020FC: begin
				q			<=			16'h8793;
		end
		32'h000020FE: begin
				q			<=			16'hFD17;
		end
		32'h00002100: begin
				q			<=			16'hB793;
		end
		32'h00002102: begin
				q			<=			16'h0017;
		end
		32'h00002104: begin
				q			<=			16'h0933;
		end
		32'h00002106: begin
				q			<=			16'h00F9;
		end
		32'h00002108: begin
				q			<=			16'h2423;
		end
		32'h0000210A: begin
				q			<=			16'h0004;
		end
		32'h0000210C: begin
				q			<=			16'h4703;
		end
		32'h0000210E: begin
				q			<=			16'h0009;
		end
		32'h00002110: begin
				q			<=			16'h0793;
		end
		32'h00002112: begin
				q			<=			16'h01F0;
		end
		32'h00002114: begin
				q			<=			16'hFE63;
		end
		32'h00002116: begin
				q			<=			16'h00E7;
		end
		32'h00002118: begin
				q			<=			16'h0A93;
		end
		32'h0000211A: begin
				q			<=			16'h0000;
		end
		32'h0000211C: begin
				q			<=			16'h0B93;
		end
		32'h0000211E: begin
				q			<=			16'h0080;
		end
		32'h00002120: begin
				q			<=			16'h0A13;
		end
		32'h00002122: begin
				q			<=			16'h02F0;
		end
		32'h00002124: begin
				q			<=			16'h0B13;
		end
		32'h00002126: begin
				q			<=			16'h02E0;
		end
		32'h00002128: begin
				q			<=			16'h0C13;
		end
		32'h0000212A: begin
				q			<=			16'h00B0;
		end
		32'h0000212C: begin
				q			<=			16'h006F;
		end
		32'h0000212E: begin
				q			<=			16'h0A00;
		end
		32'h00002130: begin
				q			<=			16'h0513;
		end
		32'h00002132: begin
				q			<=			16'h0004;
		end
		32'h00002134: begin
				q			<=			16'hF0EF;
		end
		32'h00002136: begin
				q			<=			16'hBFDF;
		end
		32'h00002138: begin
				q			<=			16'h0993;
		end
		32'h0000213A: begin
				q			<=			16'h0005;
		end
		32'h0000213C: begin
				q			<=			16'h8023;
		end
		32'h0000213E: begin
				q			<=			16'h0004;
		end
		32'h00002140: begin
				q			<=			16'h006F;
		end
		32'h00002142: begin
				q			<=			16'h1280;
		end
		32'h00002144: begin
				q			<=			16'h0513;
		end
		32'h00002146: begin
				q			<=			16'h0004;
		end
		32'h00002148: begin
				q			<=			16'hF0EF;
		end
		32'h0000214A: begin
				q			<=			16'hD51F;
		end
		32'h0000214C: begin
				q			<=			16'h1263;
		end
		32'h0000214E: begin
				q			<=			16'h0E05;
		end
		32'h00002150: begin
				q			<=			16'h5603;
		end
		32'h00002152: begin
				q			<=			16'h0004;
		end
		32'h00002154: begin
				q			<=			16'h7613;
		end
		32'h00002156: begin
				q			<=			16'h00F6;
		end
		32'h00002158: begin
				q			<=			16'h0693;
		end
		32'h0000215A: begin
				q			<=			16'h0200;
		end
		32'h0000215C: begin
				q			<=			16'h1613;
		end
		32'h0000215E: begin
				q			<=			16'h0056;
		end
		32'h00002160: begin
				q			<=			16'h2583;
		end
		32'h00002162: begin
				q			<=			16'h0104;
		end
		32'h00002164: begin
				q			<=			16'h8513;
		end
		32'h00002166: begin
				q			<=			16'h0004;
		end
		32'h00002168: begin
				q			<=			16'hF0EF;
		end
		32'h0000216A: begin
				q			<=			16'hABDF;
		end
		32'h0000216C: begin
				q			<=			16'h1663;
		end
		32'h0000216E: begin
				q			<=			16'h0C05;
		end
		32'h00002170: begin
				q			<=			16'hC783;
		end
		32'h00002172: begin
				q			<=			16'h0004;
		end
		32'h00002174: begin
				q			<=			16'h8A63;
		end
		32'h00002176: begin
				q			<=			16'h1207;
		end
		32'h00002178: begin
				q			<=			16'hC783;
		end
		32'h0000217A: begin
				q			<=			16'h00B4;
		end
		32'h0000217C: begin
				q			<=			16'hF793;
		end
		32'h0000217E: begin
				q			<=			16'h0087;
		end
		32'h00002180: begin
				q			<=			16'h92E3;
		end
		32'h00002182: begin
				q			<=			16'hFC07;
		end
		32'h00002184: begin
				q			<=			16'h2783;
		end
		32'h00002186: begin
				q			<=			16'h0044;
		end
		32'h00002188: begin
				q			<=			16'h8593;
		end
		32'h0000218A: begin
				q			<=			16'h00B7;
		end
		32'h0000218C: begin
				q			<=			16'h8713;
		end
		32'h0000218E: begin
				q			<=			16'h0004;
		end
		32'h00002190: begin
				q			<=			16'h0713;
		end
		32'h00002192: begin
				q			<=			16'h0017;
		end
		32'h00002194: begin
				q			<=			16'h8793;
		end
		32'h00002196: begin
				q			<=			16'h0017;
		end
		32'h00002198: begin
				q			<=			16'h4603;
		end
		32'h0000219A: begin
				q			<=			16'hFFF7;
		end
		32'h0000219C: begin
				q			<=			16'hC683;
		end
		32'h0000219E: begin
				q			<=			16'hFFF7;
		end
		32'h000021A0: begin
				q			<=			16'h12E3;
		end
		32'h000021A2: begin
				q			<=			16'hFAD6;
		end
		32'h000021A4: begin
				q			<=			16'h96E3;
		end
		32'h000021A6: begin
				q			<=			16'hFEF5;
		end
		32'h000021A8: begin
				q			<=			16'h2783;
		end
		32'h000021AA: begin
				q			<=			16'h0044;
		end
		32'h000021AC: begin
				q			<=			16'hC783;
		end
		32'h000021AE: begin
				q			<=			16'h00B7;
		end
		32'h000021B0: begin
				q			<=			16'h9C63;
		end
		32'h000021B2: begin
				q			<=			16'h0A07;
		end
		32'h000021B4: begin
				q			<=			16'hC783;
		end
		32'h000021B6: begin
				q			<=			16'h00B4;
		end
		32'h000021B8: begin
				q			<=			16'hF793;
		end
		32'h000021BA: begin
				q			<=			16'h0107;
		end
		32'h000021BC: begin
				q			<=			16'h8263;
		end
		32'h000021BE: begin
				q			<=			16'h0807;
		end
		32'h000021C0: begin
				q			<=			16'h8513;
		end
		32'h000021C2: begin
				q			<=			16'h0004;
		end
		32'h000021C4: begin
				q			<=			16'hF0EF;
		end
		32'h000021C6: begin
				q			<=			16'hE9DF;
		end
		32'h000021C8: begin
				q			<=			16'h2423;
		end
		32'h000021CA: begin
				q			<=			16'h00A4;
		end
		32'h000021CC: begin
				q			<=			16'h2603;
		end
		32'h000021CE: begin
				q			<=			16'h0044;
		end
		32'h000021D0: begin
				q			<=			16'h0693;
		end
		32'h000021D2: begin
				q			<=			16'h00B6;
		end
		32'h000021D4: begin
				q			<=			16'h0793;
		end
		32'h000021D6: begin
				q			<=			16'h0006;
		end
		32'h000021D8: begin
				q			<=			16'h0713;
		end
		32'h000021DA: begin
				q			<=			16'h0200;
		end
		32'h000021DC: begin
				q			<=			16'h8793;
		end
		32'h000021DE: begin
				q			<=			16'h0017;
		end
		32'h000021E0: begin
				q			<=			16'h8FA3;
		end
		32'h000021E2: begin
				q			<=			16'hFEE7;
		end
		32'h000021E4: begin
				q			<=			16'h9CE3;
		end
		32'h000021E6: begin
				q			<=			16'hFEF6;
		end
		32'h000021E8: begin
				q			<=			16'h8693;
		end
		32'h000021EA: begin
				q			<=			16'h000A;
		end
		32'h000021EC: begin
				q			<=			16'h8793;
		end
		32'h000021EE: begin
				q			<=			16'h000A;
		end
		32'h000021F0: begin
				q			<=			16'h8593;
		end
		32'h000021F2: begin
				q			<=			16'h000B;
		end
		32'h000021F4: begin
				q			<=			16'h0513;
		end
		32'h000021F6: begin
				q			<=			16'h0200;
		end
		32'h000021F8: begin
				q			<=			16'h8713;
		end
		32'h000021FA: begin
				q			<=			16'h0017;
		end
		32'h000021FC: begin
				q			<=			16'h7713;
		end
		32'h000021FE: begin
				q			<=			16'h0FF7;
		end
		32'h00002200: begin
				q			<=			16'h07B3;
		end
		32'h00002202: begin
				q			<=			16'h00F9;
		end
		32'h00002204: begin
				q			<=			16'hC783;
		end
		32'h00002206: begin
				q			<=			16'h0007;
		end
		32'h00002208: begin
				q			<=			16'h7263;
		end
		32'h0000220A: begin
				q			<=			16'h04F5;
		end
		32'h0000220C: begin
				q			<=			16'h8063;
		end
		32'h0000220E: begin
				q			<=			16'h0547;
		end
		32'h00002210: begin
				q			<=			16'h8C63;
		end
		32'h00002212: begin
				q			<=			16'h0367;
		end
		32'h00002214: begin
				q			<=			16'hFC63;
		end
		32'h00002216: begin
				q			<=			16'h02B6;
		end
		32'h00002218: begin
				q			<=			16'h8813;
		end
		32'h0000221A: begin
				q			<=			16'h0016;
		end
		32'h0000221C: begin
				q			<=			16'h06B3;
		end
		32'h0000221E: begin
				q			<=			16'h00D6;
		end
		32'h00002220: begin
				q			<=			16'h8023;
		end
		32'h00002222: begin
				q			<=			16'h00F6;
		end
		32'h00002224: begin
				q			<=			16'h7693;
		end
		32'h00002226: begin
				q			<=			16'h0FF8;
		end
		32'h00002228: begin
				q			<=			16'h0793;
		end
		32'h0000222A: begin
				q			<=			16'h0007;
		end
		32'h0000222C: begin
				q			<=			16'hF06F;
		end
		32'h0000222E: begin
				q			<=			16'hFCDF;
		end
		32'h00002230: begin
				q			<=			16'h0993;
		end
		32'h00002232: begin
				q			<=			16'h0005;
		end
		32'h00002234: begin
				q			<=			16'h006F;
		end
		32'h00002236: begin
				q			<=			16'h0340;
		end
		32'h00002238: begin
				q			<=			16'h0993;
		end
		32'h0000223A: begin
				q			<=			16'h0010;
		end
		32'h0000223C: begin
				q			<=			16'h006F;
		end
		32'h0000223E: begin
				q			<=			16'h02C0;
		end
		32'h00002240: begin
				q			<=			16'h0993;
		end
		32'h00002242: begin
				q			<=			16'h0030;
		end
		32'h00002244: begin
				q			<=			16'h006F;
		end
		32'h00002246: begin
				q			<=			16'h0240;
		end
		32'h00002248: begin
				q			<=			16'h8A63;
		end
		32'h0000224A: begin
				q			<=			16'h0575;
		end
		32'h0000224C: begin
				q			<=			16'h0933;
		end
		32'h0000224E: begin
				q			<=			16'h00E9;
		end
		32'h00002250: begin
				q			<=			16'hB793;
		end
		32'h00002252: begin
				q			<=			16'h0217;
		end
		32'h00002254: begin
				q			<=			16'h05A3;
		end
		32'h00002256: begin
				q			<=			16'h00F6;
		end
		32'h00002258: begin
				q			<=			16'h0513;
		end
		32'h0000225A: begin
				q			<=			16'h0004;
		end
		32'h0000225C: begin
				q			<=			16'hF0EF;
		end
		32'h0000225E: begin
				q			<=			16'hAD5F;
		end
		32'h00002260: begin
				q			<=			16'h0993;
		end
		32'h00002262: begin
				q			<=			16'h0005;
		end
		32'h00002264: begin
				q			<=			16'h06E3;
		end
		32'h00002266: begin
				q			<=			16'hEE05;
		end
		32'h00002268: begin
				q			<=			16'h8513;
		end
		32'h0000226A: begin
				q			<=			16'h0009;
		end
		32'h0000226C: begin
				q			<=			16'h2083;
		end
		32'h0000226E: begin
				q			<=			16'h02C1;
		end
		32'h00002270: begin
				q			<=			16'h2403;
		end
		32'h00002272: begin
				q			<=			16'h0281;
		end
		32'h00002274: begin
				q			<=			16'h2483;
		end
		32'h00002276: begin
				q			<=			16'h0241;
		end
		32'h00002278: begin
				q			<=			16'h2903;
		end
		32'h0000227A: begin
				q			<=			16'h0201;
		end
		32'h0000227C: begin
				q			<=			16'h2983;
		end
		32'h0000227E: begin
				q			<=			16'h01C1;
		end
		32'h00002280: begin
				q			<=			16'h2A03;
		end
		32'h00002282: begin
				q			<=			16'h0181;
		end
		32'h00002284: begin
				q			<=			16'h2A83;
		end
		32'h00002286: begin
				q			<=			16'h0141;
		end
		32'h00002288: begin
				q			<=			16'h2B03;
		end
		32'h0000228A: begin
				q			<=			16'h0101;
		end
		32'h0000228C: begin
				q			<=			16'h2B83;
		end
		32'h0000228E: begin
				q			<=			16'h00C1;
		end
		32'h00002290: begin
				q			<=			16'h2C03;
		end
		32'h00002292: begin
				q			<=			16'h0081;
		end
		32'h00002294: begin
				q			<=			16'h0113;
		end
		32'h00002296: begin
				q			<=			16'h0301;
		end
		32'h00002298: begin
				q			<=			16'h8067;
		end
		32'h0000229A: begin
				q			<=			16'h0000;
		end
		32'h0000229C: begin
				q			<=			16'h8693;
		end
		32'h0000229E: begin
				q			<=			16'h0005;
		end
		32'h000022A0: begin
				q			<=			16'h0593;
		end
		32'h000022A2: begin
				q			<=			16'h000C;
		end
		32'h000022A4: begin
				q			<=			16'hF06F;
		end
		32'h000022A6: begin
				q			<=			16'hF85F;
		end
		32'h000022A8: begin
				q			<=			16'h0993;
		end
		32'h000022AA: begin
				q			<=			16'h0030;
		end
		32'h000022AC: begin
				q			<=			16'hF06F;
		end
		32'h000022AE: begin
				q			<=			16'hFBDF;
		end
		32'h000022B0: begin
				q			<=			16'h0000;
		end
		32'h000022B2: begin
				q			<=			16'h0000;
		end
		32'h000022B4: begin
				q			<=			16'h0113;
		end
		32'h000022B6: begin
				q			<=			16'hFB01;
		end
		32'h000022B8: begin
				q			<=			16'h2623;
		end
		32'h000022BA: begin
				q			<=			16'h0411;
		end
		32'h000022BC: begin
				q			<=			16'h2423;
		end
		32'h000022BE: begin
				q			<=			16'h0481;
		end
		32'h000022C0: begin
				q			<=			16'h2223;
		end
		32'h000022C2: begin
				q			<=			16'h0491;
		end
		32'h000022C4: begin
				q			<=			16'h2023;
		end
		32'h000022C6: begin
				q			<=			16'h0521;
		end
		32'h000022C8: begin
				q			<=			16'h2E23;
		end
		32'h000022CA: begin
				q			<=			16'h0331;
		end
		32'h000022CC: begin
				q			<=			16'h2C23;
		end
		32'h000022CE: begin
				q			<=			16'h0341;
		end
		32'h000022D0: begin
				q			<=			16'h2A23;
		end
		32'h000022D2: begin
				q			<=			16'h0351;
		end
		32'h000022D4: begin
				q			<=			16'h0413;
		end
		32'h000022D6: begin
				q			<=			16'h0005;
		end
		32'h000022D8: begin
				q			<=			16'h17B7;
		end
		32'h000022DA: begin
				q			<=			16'h0001;
		end
		32'h000022DC: begin
				q			<=			16'hAE23;
		end
		32'h000022DE: begin
				q			<=			16'hF807;
		end
		32'h000022E0: begin
				q			<=			16'hF0EF;
		end
		32'h000022E2: begin
				q			<=			16'h939F;
		end
		32'h000022E4: begin
				q			<=			16'h7513;
		end
		32'h000022E6: begin
				q			<=			16'h0015;
		end
		32'h000022E8: begin
				q			<=			16'h0793;
		end
		32'h000022EA: begin
				q			<=			16'h0020;
		end
		32'h000022EC: begin
				q			<=			16'h1663;
		end
		32'h000022EE: begin
				q			<=			16'h1205;
		end
		32'h000022F0: begin
				q			<=			16'h0593;
		end
		32'h000022F2: begin
				q			<=			16'h0000;
		end
		32'h000022F4: begin
				q			<=			16'h0513;
		end
		32'h000022F6: begin
				q			<=			16'h00C1;
		end
		32'h000022F8: begin
				q			<=			16'hF0EF;
		end
		32'h000022FA: begin
				q			<=			16'hC71F;
		end
		32'h000022FC: begin
				q			<=			16'h0793;
		end
		32'h000022FE: begin
				q			<=			16'h0010;
		end
		32'h00002300: begin
				q			<=			16'h0493;
		end
		32'h00002302: begin
				q			<=			16'h0000;
		end
		32'h00002304: begin
				q			<=			16'h0E63;
		end
		32'h00002306: begin
				q			<=			16'h12F5;
		end
		32'h00002308: begin
				q			<=			16'h0713;
		end
		32'h0000230A: begin
				q			<=			16'h0030;
		end
		32'h0000230C: begin
				q			<=			16'h0793;
		end
		32'h0000230E: begin
				q			<=			16'h0010;
		end
		32'h00002310: begin
				q			<=			16'h0463;
		end
		32'h00002312: begin
				q			<=			16'h10E5;
		end
		32'h00002314: begin
				q			<=			16'h0793;
		end
		32'h00002316: begin
				q			<=			16'h0060;
		end
		32'h00002318: begin
				q			<=			16'h1063;
		end
		32'h0000231A: begin
				q			<=			16'h1005;
		end
		32'h0000231C: begin
				q			<=			16'h0693;
		end
		32'h0000231E: begin
				q			<=			16'h0240;
		end
		32'h00002320: begin
				q			<=			16'h0613;
		end
		32'h00002322: begin
				q			<=			16'h00D0;
		end
		32'h00002324: begin
				q			<=			16'h8593;
		end
		32'h00002326: begin
				q			<=			16'h0004;
		end
		32'h00002328: begin
				q			<=			16'h0513;
		end
		32'h0000232A: begin
				q			<=			16'h00C1;
		end
		32'h0000232C: begin
				q			<=			16'hF0EF;
		end
		32'h0000232E: begin
				q			<=			16'h8F9F;
		end
		32'h00002330: begin
				q			<=			16'h0793;
		end
		32'h00002332: begin
				q			<=			16'h0010;
		end
		32'h00002334: begin
				q			<=			16'h1263;
		end
		32'h00002336: begin
				q			<=			16'h0E05;
		end
		32'h00002338: begin
				q			<=			16'h4503;
		end
		32'h0000233A: begin
				q			<=			16'h0161;
		end
		32'h0000233C: begin
				q			<=			16'h1513;
		end
		32'h0000233E: begin
				q			<=			16'h0085;
		end
		32'h00002340: begin
				q			<=			16'h4783;
		end
		32'h00002342: begin
				q			<=			16'h0151;
		end
		32'h00002344: begin
				q			<=			16'h6533;
		end
		32'h00002346: begin
				q			<=			16'h00F5;
		end
		32'h00002348: begin
				q			<=			16'h1663;
		end
		32'h0000234A: begin
				q			<=			16'h0005;
		end
		32'h0000234C: begin
				q			<=			16'h0513;
		end
		32'h0000234E: begin
				q			<=			16'h0231;
		end
		32'h00002350: begin
				q			<=			16'hF0EF;
		end
		32'h00002352: begin
				q			<=			16'h979F;
		end
		32'h00002354: begin
				q			<=			16'h4983;
		end
		32'h00002356: begin
				q			<=			16'h00F1;
		end
		32'h00002358: begin
				q			<=			16'h89B3;
		end
		32'h0000235A: begin
				q			<=			16'h02A9;
		end
		32'h0000235C: begin
				q			<=			16'h4783;
		end
		32'h0000235E: begin
				q			<=			16'h00E1;
		end
		32'h00002360: begin
				q			<=			16'h9793;
		end
		32'h00002362: begin
				q			<=			16'h0087;
		end
		32'h00002364: begin
				q			<=			16'h4A83;
		end
		32'h00002366: begin
				q			<=			16'h00D1;
		end
		32'h00002368: begin
				q			<=			16'hEAB3;
		end
		32'h0000236A: begin
				q			<=			16'h0157;
		end
		32'h0000236C: begin
				q			<=			16'h84B3;
		end
		32'h0000236E: begin
				q			<=			16'h009A;
		end
		32'h00002370: begin
				q			<=			16'h2623;
		end
		32'h00002372: begin
				q			<=			16'h0094;
		end
		32'h00002374: begin
				q			<=			16'h4A03;
		end
		32'h00002376: begin
				q			<=			16'h00C1;
		end
		32'h00002378: begin
				q			<=			16'h0123;
		end
		32'h0000237A: begin
				q			<=			16'h0144;
		end
		32'h0000237C: begin
				q			<=			16'h4903;
		end
		32'h0000237E: begin
				q			<=			16'h0111;
		end
		32'h00002380: begin
				q			<=			16'h1913;
		end
		32'h00002382: begin
				q			<=			16'h0089;
		end
		32'h00002384: begin
				q			<=			16'h4783;
		end
		32'h00002386: begin
				q			<=			16'h0101;
		end
		32'h00002388: begin
				q			<=			16'h6933;
		end
		32'h0000238A: begin
				q			<=			16'h00F9;
		end
		32'h0000238C: begin
				q			<=			16'h1223;
		end
		32'h0000238E: begin
				q			<=			16'h0124;
		end
		32'h00002390: begin
				q			<=			16'h4503;
		end
		32'h00002392: begin
				q			<=			16'h0131;
		end
		32'h00002394: begin
				q			<=			16'h1513;
		end
		32'h00002396: begin
				q			<=			16'h0085;
		end
		32'h00002398: begin
				q			<=			16'h4783;
		end
		32'h0000239A: begin
				q			<=			16'h0121;
		end
		32'h0000239C: begin
				q			<=			16'h6533;
		end
		32'h0000239E: begin
				q			<=			16'h00F5;
		end
		32'h000023A0: begin
				q			<=			16'h1663;
		end
		32'h000023A2: begin
				q			<=			16'h0005;
		end
		32'h000023A4: begin
				q			<=			16'h0513;
		end
		32'h000023A6: begin
				q			<=			16'h01F1;
		end
		32'h000023A8: begin
				q			<=			16'hF0EF;
		end
		32'h000023AA: begin
				q			<=			16'h921F;
		end
		32'h000023AC: begin
				q			<=			16'h5913;
		end
		32'h000023AE: begin
				q			<=			16'h0049;
		end
		32'h000023B0: begin
				q			<=			16'h07B3;
		end
		32'h000023B2: begin
				q			<=			16'h4155;
		end
		32'h000023B4: begin
				q			<=			16'h87B3;
		end
		32'h000023B6: begin
				q			<=			16'h4137;
		end
		32'h000023B8: begin
				q			<=			16'h87B3;
		end
		32'h000023BA: begin
				q			<=			16'h4127;
		end
		32'h000023BC: begin
				q			<=			16'hD7B3;
		end
		32'h000023BE: begin
				q			<=			16'h0347;
		end
		32'h000023C0: begin
				q			<=			16'h8693;
		end
		32'h000023C2: begin
				q			<=			16'h0027;
		end
		32'h000023C4: begin
				q			<=			16'h2423;
		end
		32'h000023C6: begin
				q			<=			16'h00D4;
		end
		32'h000023C8: begin
				q			<=			16'hF737;
		end
		32'h000023CA: begin
				q			<=			16'hFFFF;
		end
		32'h000023CC: begin
				q			<=			16'h0713;
		end
		32'h000023CE: begin
				q			<=			16'h00A7;
		end
		32'h000023D0: begin
				q			<=			16'h87B3;
		end
		32'h000023D2: begin
				q			<=			16'h00E7;
		end
		32'h000023D4: begin
				q			<=			16'hF737;
		end
		32'h000023D6: begin
				q			<=			16'h0000;
		end
		32'h000023D8: begin
				q			<=			16'h0713;
		end
		32'h000023DA: begin
				q			<=			16'hFFE7;
		end
		32'h000023DC: begin
				q			<=			16'h6463;
		end
		32'h000023DE: begin
				q			<=			16'h0AF7;
		end
		32'h000023E0: begin
				q			<=			16'h07B7;
		end
		32'h000023E2: begin
				q			<=			16'h0001;
		end
		32'h000023E4: begin
				q			<=			16'h8793;
		end
		32'h000023E6: begin
				q			<=			16'hFF67;
		end
		32'h000023E8: begin
				q			<=			16'hE463;
		end
		32'h000023EA: begin
				q			<=			16'h0CD7;
		end
		32'h000023EC: begin
				q			<=			16'h0793;
		end
		32'h000023EE: begin
				q			<=			16'h0020;
		end
		32'h000023F0: begin
				q			<=			16'h0023;
		end
		32'h000023F2: begin
				q			<=			16'h00F4;
		end
		32'h000023F4: begin
				q			<=			16'h87B3;
		end
		32'h000023F6: begin
				q			<=			16'h0134;
		end
		32'h000023F8: begin
				q			<=			16'h2823;
		end
		32'h000023FA: begin
				q			<=			16'h00F4;
		end
		32'h000023FC: begin
				q			<=			16'h84B3;
		end
		32'h000023FE: begin
				q			<=			16'h0124;
		end
		32'h00002400: begin
				q			<=			16'h8533;
		end
		32'h00002402: begin
				q			<=			16'h0134;
		end
		32'h00002404: begin
				q			<=			16'h2A23;
		end
		32'h00002406: begin
				q			<=			16'h00A4;
		end
		32'h00002408: begin
				q			<=			16'h00A3;
		end
		32'h0000240A: begin
				q			<=			16'h0004;
		end
		32'h0000240C: begin
				q			<=			16'h17B7;
		end
		32'h0000240E: begin
				q			<=			16'h0001;
		end
		32'h00002410: begin
				q			<=			16'hAE23;
		end
		32'h00002412: begin
				q			<=			16'hF887;
		end
		32'h00002414: begin
				q			<=			16'h0793;
		end
		32'h00002416: begin
				q			<=			16'h0000;
		end
		32'h00002418: begin
				q			<=			16'h8513;
		end
		32'h0000241A: begin
				q			<=			16'h0007;
		end
		32'h0000241C: begin
				q			<=			16'h2083;
		end
		32'h0000241E: begin
				q			<=			16'h04C1;
		end
		32'h00002420: begin
				q			<=			16'h2403;
		end
		32'h00002422: begin
				q			<=			16'h0481;
		end
		32'h00002424: begin
				q			<=			16'h2483;
		end
		32'h00002426: begin
				q			<=			16'h0441;
		end
		32'h00002428: begin
				q			<=			16'h2903;
		end
		32'h0000242A: begin
				q			<=			16'h0401;
		end
		32'h0000242C: begin
				q			<=			16'h2983;
		end
		32'h0000242E: begin
				q			<=			16'h03C1;
		end
		32'h00002430: begin
				q			<=			16'h2A03;
		end
		32'h00002432: begin
				q			<=			16'h0381;
		end
		32'h00002434: begin
				q			<=			16'h2A83;
		end
		32'h00002436: begin
				q			<=			16'h0341;
		end
		32'h00002438: begin
				q			<=			16'h0113;
		end
		32'h0000243A: begin
				q			<=			16'h0501;
		end
		32'h0000243C: begin
				q			<=			16'h8067;
		end
		32'h0000243E: begin
				q			<=			16'h0000;
		end
		32'h00002440: begin
				q			<=			16'h0693;
		end
		32'h00002442: begin
				q			<=			16'h0100;
		end
		32'h00002444: begin
				q			<=			16'h0613;
		end
		32'h00002446: begin
				q			<=			16'h1BE0;
		end
		32'h00002448: begin
				q			<=			16'h0593;
		end
		32'h0000244A: begin
				q			<=			16'h0000;
		end
		32'h0000244C: begin
				q			<=			16'h0513;
		end
		32'h0000244E: begin
				q			<=			16'h00C1;
		end
		32'h00002450: begin
				q			<=			16'hF0EF;
		end
		32'h00002452: begin
				q			<=			16'hFD4F;
		end
		32'h00002454: begin
				q			<=			16'h0793;
		end
		32'h00002456: begin
				q			<=			16'h0010;
		end
		32'h00002458: begin
				q			<=			16'h10E3;
		end
		32'h0000245A: begin
				q			<=			16'hFC05;
		end
		32'h0000245C: begin
				q			<=			16'h4703;
		end
		32'h0000245E: begin
				q			<=			16'h0101;
		end
		32'h00002460: begin
				q			<=			16'h0793;
		end
		32'h00002462: begin
				q			<=			16'h0060;
		end
		32'h00002464: begin
				q			<=			16'h0AE3;
		end
		32'h00002466: begin
				q			<=			16'hFA07;
		end
		32'h00002468: begin
				q			<=			16'h0513;
		end
		32'h0000246A: begin
				q			<=			16'h0141;
		end
		32'h0000246C: begin
				q			<=			16'hF0EF;
		end
		32'h0000246E: begin
				q			<=			16'h85DF;
		end
		32'h00002470: begin
				q			<=			16'h0493;
		end
		32'h00002472: begin
				q			<=			16'h0005;
		end
		32'h00002474: begin
				q			<=			16'h0593;
		end
		32'h00002476: begin
				q			<=			16'h0005;
		end
		32'h00002478: begin
				q			<=			16'h0513;
		end
		32'h0000247A: begin
				q			<=			16'h00C1;
		end
		32'h0000247C: begin
				q			<=			16'hF0EF;
		end
		32'h0000247E: begin
				q			<=			16'hAEDF;
		end
		32'h00002480: begin
				q			<=			16'hF06F;
		end
		32'h00002482: begin
				q			<=			16'hE89F;
		end
		32'h00002484: begin
				q			<=			16'h07B7;
		end
		32'h00002486: begin
				q			<=			16'h0001;
		end
		32'h00002488: begin
				q			<=			16'h8793;
		end
		32'h0000248A: begin
				q			<=			16'hFF67;
		end
		32'h0000248C: begin
				q			<=			16'hFE63;
		end
		32'h0000248E: begin
				q			<=			16'h00D7;
		end
		32'h00002490: begin
				q			<=			16'h0793;
		end
		32'h00002492: begin
				q			<=			16'h0030;
		end
		32'h00002494: begin
				q			<=			16'h0023;
		end
		32'h00002496: begin
				q			<=			16'h00F4;
		end
		32'h00002498: begin
				q			<=			16'h0513;
		end
		32'h0000249A: begin
				q			<=			16'h02B1;
		end
		32'h0000249C: begin
				q			<=			16'hF0EF;
		end
		32'h0000249E: begin
				q			<=			16'h82DF;
		end
		32'h000024A0: begin
				q			<=			16'h2823;
		end
		32'h000024A2: begin
				q			<=			16'h00A4;
		end
		32'h000024A4: begin
				q			<=			16'hF06F;
		end
		32'h000024A6: begin
				q			<=			16'hF59F;
		end
		32'h000024A8: begin
				q			<=			16'h0793;
		end
		32'h000024AA: begin
				q			<=			16'h0060;
		end
		32'h000024AC: begin
				q			<=			16'hF06F;
		end
		32'h000024AE: begin
				q			<=			16'hF6DF;
		end
		32'h000024B0: begin
				q			<=			16'h0793;
		end
		32'h000024B2: begin
				q			<=			16'h0030;
		end
		32'h000024B4: begin
				q			<=			16'h0023;
		end
		32'h000024B6: begin
				q			<=			16'h00F4;
		end
		32'h000024B8: begin
				q			<=			16'hF06F;
		end
		32'h000024BA: begin
				q			<=			16'hFE1F;
		end
		32'h000024BC: begin
				q			<=			16'h0000;
		end
		32'h000024BE: begin
				q			<=			16'h0000;
		end
		32'h000024C0: begin
				q			<=			16'h0113;
		end
		32'h000024C2: begin
				q			<=			16'hFB01;
		end
		32'h000024C4: begin
				q			<=			16'h2623;
		end
		32'h000024C6: begin
				q			<=			16'h0411;
		end
		32'h000024C8: begin
				q			<=			16'h2423;
		end
		32'h000024CA: begin
				q			<=			16'h0481;
		end
		32'h000024CC: begin
				q			<=			16'h2223;
		end
		32'h000024CE: begin
				q			<=			16'h0491;
		end
		32'h000024D0: begin
				q			<=			16'h17B7;
		end
		32'h000024D2: begin
				q			<=			16'h0001;
		end
		32'h000024D4: begin
				q			<=			16'hA403;
		end
		32'h000024D6: begin
				q			<=			16'hF9C7;
		end
		32'h000024D8: begin
				q			<=			16'h0493;
		end
		32'h000024DA: begin
				q			<=			16'h0050;
		end
		32'h000024DC: begin
				q			<=			16'h0063;
		end
		32'h000024DE: begin
				q			<=			16'h0604;
		end
		32'h000024E0: begin
				q			<=			16'h0613;
		end
		32'h000024E2: begin
				q			<=			16'h0005;
		end
		32'h000024E4: begin
				q			<=			16'h00A3;
		end
		32'h000024E6: begin
				q			<=			16'h0004;
		end
		32'h000024E8: begin
				q			<=			16'h0793;
		end
		32'h000024EA: begin
				q			<=			16'h0201;
		end
		32'h000024EC: begin
				q			<=			16'h2823;
		end
		32'h000024EE: begin
				q			<=			16'h02F1;
		end
		32'h000024F0: begin
				q			<=			16'h0593;
		end
		32'h000024F2: begin
				q			<=			16'h0001;
		end
		32'h000024F4: begin
				q			<=			16'h0513;
		end
		32'h000024F6: begin
				q			<=			16'h02C1;
		end
		32'h000024F8: begin
				q			<=			16'hF0EF;
		end
		32'h000024FA: begin
				q			<=			16'hBB5F;
		end
		32'h000024FC: begin
				q			<=			16'h0493;
		end
		32'h000024FE: begin
				q			<=			16'h0005;
		end
		32'h00002500: begin
				q			<=			16'h1E63;
		end
		32'h00002502: begin
				q			<=			16'h0205;
		end
		32'h00002504: begin
				q			<=			16'h4783;
		end
		32'h00002506: begin
				q			<=			16'h0001;
		end
		32'h00002508: begin
				q			<=			16'h8663;
		end
		32'h0000250A: begin
				q			<=			16'h0407;
		end
		32'h0000250C: begin
				q			<=			16'h4783;
		end
		32'h0000250E: begin
				q			<=			16'h00B1;
		end
		32'h00002510: begin
				q			<=			16'hF793;
		end
		32'h00002512: begin
				q			<=			16'h0107;
		end
		32'h00002514: begin
				q			<=			16'h9463;
		end
		32'h00002516: begin
				q			<=			16'h0407;
		end
		32'h00002518: begin
				q			<=			16'h0513;
		end
		32'h0000251A: begin
				q			<=			16'h0001;
		end
		32'h0000251C: begin
				q			<=			16'hF0EF;
		end
		32'h0000251E: begin
				q			<=			16'hB45F;
		end
		32'h00002520: begin
				q			<=			16'h2023;
		end
		32'h00002522: begin
				q			<=			16'h02A4;
		end
		32'h00002524: begin
				q			<=			16'h0513;
		end
		32'h00002526: begin
				q			<=			16'h01C1;
		end
		32'h00002528: begin
				q			<=			16'hF0EF;
		end
		32'h0000252A: begin
				q			<=			16'hFA0F;
		end
		32'h0000252C: begin
				q			<=			16'h2E23;
		end
		32'h0000252E: begin
				q			<=			16'h00A4;
		end
		32'h00002530: begin
				q			<=			16'h2C23;
		end
		32'h00002532: begin
				q			<=			16'h0004;
		end
		32'h00002534: begin
				q			<=			16'h0793;
		end
		32'h00002536: begin
				q			<=			16'h0010;
		end
		32'h00002538: begin
				q			<=			16'h00A3;
		end
		32'h0000253A: begin
				q			<=			16'h00F4;
		end
		32'h0000253C: begin
				q			<=			16'h8513;
		end
		32'h0000253E: begin
				q			<=			16'h0004;
		end
		32'h00002540: begin
				q			<=			16'h2083;
		end
		32'h00002542: begin
				q			<=			16'h04C1;
		end
		32'h00002544: begin
				q			<=			16'h2403;
		end
		32'h00002546: begin
				q			<=			16'h0481;
		end
		32'h00002548: begin
				q			<=			16'h2483;
		end
		32'h0000254A: begin
				q			<=			16'h0441;
		end
		32'h0000254C: begin
				q			<=			16'h0113;
		end
		32'h0000254E: begin
				q			<=			16'h0501;
		end
		32'h00002550: begin
				q			<=			16'h8067;
		end
		32'h00002552: begin
				q			<=			16'h0000;
		end
		32'h00002554: begin
				q			<=			16'h0493;
		end
		32'h00002556: begin
				q			<=			16'h0030;
		end
		32'h00002558: begin
				q			<=			16'hF06F;
		end
		32'h0000255A: begin
				q			<=			16'hFE5F;
		end
		32'h0000255C: begin
				q			<=			16'h0493;
		end
		32'h0000255E: begin
				q			<=			16'h0030;
		end
		32'h00002560: begin
				q			<=			16'hF06F;
		end
		32'h00002562: begin
				q			<=			16'hFDDF;
		end
		32'h00002564: begin
				q			<=			16'h0000;
		end
		32'h00002566: begin
				q			<=			16'h0000;
		end
		32'h00002568: begin
				q			<=			16'h0113;
		end
		32'h0000256A: begin
				q			<=			16'hFE01;
		end
		32'h0000256C: begin
				q			<=			16'h2E23;
		end
		32'h0000256E: begin
				q			<=			16'h0011;
		end
		32'h00002570: begin
				q			<=			16'h2C23;
		end
		32'h00002572: begin
				q			<=			16'h0081;
		end
		32'h00002574: begin
				q			<=			16'h2A23;
		end
		32'h00002576: begin
				q			<=			16'h0091;
		end
		32'h00002578: begin
				q			<=			16'h2823;
		end
		32'h0000257A: begin
				q			<=			16'h0121;
		end
		32'h0000257C: begin
				q			<=			16'h2623;
		end
		32'h0000257E: begin
				q			<=			16'h0131;
		end
		32'h00002580: begin
				q			<=			16'h2423;
		end
		32'h00002582: begin
				q			<=			16'h0141;
		end
		32'h00002584: begin
				q			<=			16'h2223;
		end
		32'h00002586: begin
				q			<=			16'h0151;
		end
		32'h00002588: begin
				q			<=			16'h2023;
		end
		32'h0000258A: begin
				q			<=			16'h0161;
		end
		32'h0000258C: begin
				q			<=			16'h17B7;
		end
		32'h0000258E: begin
				q			<=			16'h0001;
		end
		32'h00002590: begin
				q			<=			16'hA403;
		end
		32'h00002592: begin
				q			<=			16'hF9C7;
		end
		32'h00002594: begin
				q			<=			16'h2023;
		end
		32'h00002596: begin
				q			<=			16'h0006;
		end
		32'h00002598: begin
				q			<=			16'h0A63;
		end
		32'h0000259A: begin
				q			<=			16'h1204;
		end
		32'h0000259C: begin
				q			<=			16'h0993;
		end
		32'h0000259E: begin
				q			<=			16'h0005;
		end
		32'h000025A0: begin
				q			<=			16'h0A13;
		end
		32'h000025A2: begin
				q			<=			16'h0006;
		end
		32'h000025A4: begin
				q			<=			16'h4783;
		end
		32'h000025A6: begin
				q			<=			16'h0014;
		end
		32'h000025A8: begin
				q			<=			16'hF793;
		end
		32'h000025AA: begin
				q			<=			16'h0017;
		end
		32'h000025AC: begin
				q			<=			16'h0513;
		end
		32'h000025AE: begin
				q			<=			16'h0040;
		end
		32'h000025B0: begin
				q			<=			16'h8663;
		end
		32'h000025B2: begin
				q			<=			16'h0E07;
		end
		32'h000025B4: begin
				q			<=			16'h2903;
		end
		32'h000025B6: begin
				q			<=			16'h01C4;
		end
		32'h000025B8: begin
				q			<=			16'h2783;
		end
		32'h000025BA: begin
				q			<=			16'h0184;
		end
		32'h000025BC: begin
				q			<=			16'h0933;
		end
		32'h000025BE: begin
				q			<=			16'h40F9;
		end
		32'h000025C0: begin
				q			<=			16'hF463;
		end
		32'h000025C2: begin
				q			<=			16'h0125;
		end
		32'h000025C4: begin
				q			<=			16'h8913;
		end
		32'h000025C6: begin
				q			<=			16'h0005;
		end
		32'h000025C8: begin
				q			<=			16'h0663;
		end
		32'h000025CA: begin
				q			<=			16'h1009;
		end
		32'h000025CC: begin
				q			<=			16'h0B13;
		end
		32'h000025CE: begin
				q			<=			16'h0010;
		end
		32'h000025D0: begin
				q			<=			16'h0A93;
		end
		32'h000025D2: begin
				q			<=			16'h2000;
		end
		32'h000025D4: begin
				q			<=			16'h006F;
		end
		32'h000025D6: begin
				q			<=			16'h0780;
		end
		32'h000025D8: begin
				q			<=			16'h2503;
		end
		32'h000025DA: begin
				q			<=			16'h0244;
		end
		32'h000025DC: begin
				q			<=			16'hF0EF;
		end
		32'h000025DE: begin
				q			<=			16'hFE4F;
		end
		32'h000025E0: begin
				q			<=			16'h7E63;
		end
		32'h000025E2: begin
				q			<=			16'h08AB;
		end
		32'h000025E4: begin
				q			<=			16'h2223;
		end
		32'h000025E6: begin
				q			<=			16'h02A4;
		end
		32'h000025E8: begin
				q			<=			16'h2503;
		end
		32'h000025EA: begin
				q			<=			16'h0244;
		end
		32'h000025EC: begin
				q			<=			16'hF0EF;
		end
		32'h000025EE: begin
				q			<=			16'hF0CF;
		end
		32'h000025F0: begin
				q			<=			16'h0C63;
		end
		32'h000025F2: begin
				q			<=			16'h0805;
		end
		32'h000025F4: begin
				q			<=			16'h84B3;
		end
		32'h000025F6: begin
				q			<=			16'h00A4;
		end
		32'h000025F8: begin
				q			<=			16'h2423;
		end
		32'h000025FA: begin
				q			<=			16'h0294;
		end
		32'h000025FC: begin
				q			<=			16'h2603;
		end
		32'h000025FE: begin
				q			<=			16'h0184;
		end
		32'h00002600: begin
				q			<=			16'h7613;
		end
		32'h00002602: begin
				q			<=			16'h1FF6;
		end
		32'h00002604: begin
				q			<=			16'h84B3;
		end
		32'h00002606: begin
				q			<=			16'h40CA;
		end
		32'h00002608: begin
				q			<=			16'h7463;
		end
		32'h0000260A: begin
				q			<=			16'h0099;
		end
		32'h0000260C: begin
				q			<=			16'h0493;
		end
		32'h0000260E: begin
				q			<=			16'h0009;
		end
		32'h00002610: begin
				q			<=			16'h8693;
		end
		32'h00002612: begin
				q			<=			16'h0004;
		end
		32'h00002614: begin
				q			<=			16'h2583;
		end
		32'h00002616: begin
				q			<=			16'h0284;
		end
		32'h00002618: begin
				q			<=			16'h8513;
		end
		32'h0000261A: begin
				q			<=			16'h0009;
		end
		32'h0000261C: begin
				q			<=			16'hF0EF;
		end
		32'h0000261E: begin
				q			<=			16'hE08F;
		end
		32'h00002620: begin
				q			<=			16'h1A63;
		end
		32'h00002622: begin
				q			<=			16'h0605;
		end
		32'h00002624: begin
				q			<=			16'h2783;
		end
		32'h00002626: begin
				q			<=			16'h0184;
		end
		32'h00002628: begin
				q			<=			16'h87B3;
		end
		32'h0000262A: begin
				q			<=			16'h0097;
		end
		32'h0000262C: begin
				q			<=			16'h2C23;
		end
		32'h0000262E: begin
				q			<=			16'h00F4;
		end
		32'h00002630: begin
				q			<=			16'h0933;
		end
		32'h00002632: begin
				q			<=			16'h4099;
		end
		32'h00002634: begin
				q			<=			16'h2783;
		end
		32'h00002636: begin
				q			<=			16'h000A;
		end
		32'h00002638: begin
				q			<=			16'h87B3;
		end
		32'h0000263A: begin
				q			<=			16'h0097;
		end
		32'h0000263C: begin
				q			<=			16'h2023;
		end
		32'h0000263E: begin
				q			<=			16'h00FA;
		end
		32'h00002640: begin
				q			<=			16'h8463;
		end
		32'h00002642: begin
				q			<=			16'h0009;
		end
		32'h00002644: begin
				q			<=			16'h89B3;
		end
		32'h00002646: begin
				q			<=			16'h0099;
		end
		32'h00002648: begin
				q			<=			16'h0E63;
		end
		32'h0000264A: begin
				q			<=			16'h0609;
		end
		32'h0000264C: begin
				q			<=			16'h2783;
		end
		32'h0000264E: begin
				q			<=			16'h0184;
		end
		32'h00002650: begin
				q			<=			16'hF713;
		end
		32'h00002652: begin
				q			<=			16'h1FF7;
		end
		32'h00002654: begin
				q			<=			16'h14E3;
		end
		32'h00002656: begin
				q			<=			16'hFA07;
		end
		32'h00002658: begin
				q			<=			16'h4483;
		end
		32'h0000265A: begin
				q			<=			16'h0024;
		end
		32'h0000265C: begin
				q			<=			16'h8493;
		end
		32'h0000265E: begin
				q			<=			16'hFFF4;
		end
		32'h00002660: begin
				q			<=			16'hD513;
		end
		32'h00002662: begin
				q			<=			16'h0097;
		end
		32'h00002664: begin
				q			<=			16'hF4B3;
		end
		32'h00002666: begin
				q			<=			16'h00A4;
		end
		32'h00002668: begin
				q			<=			16'hF493;
		end
		32'h0000266A: begin
				q			<=			16'h0FF4;
		end
		32'h0000266C: begin
				q			<=			16'h9EE3;
		end
		32'h0000266E: begin
				q			<=			16'hF604;
		end
		32'h00002670: begin
				q			<=			16'h94E3;
		end
		32'h00002672: begin
				q			<=			16'hF607;
		end
		32'h00002674: begin
				q			<=			16'h2503;
		end
		32'h00002676: begin
				q			<=			16'h0204;
		end
		32'h00002678: begin
				q			<=			16'hF06F;
		end
		32'h0000267A: begin
				q			<=			16'hF69F;
		end
		32'h0000267C: begin
				q			<=			16'h00A3;
		end
		32'h0000267E: begin
				q			<=			16'h0004;
		end
		32'h00002680: begin
				q			<=			16'h0513;
		end
		32'h00002682: begin
				q			<=			16'h0010;
		end
		32'h00002684: begin
				q			<=			16'h006F;
		end
		32'h00002686: begin
				q			<=			16'h0180;
		end
		32'h00002688: begin
				q			<=			16'h00A3;
		end
		32'h0000268A: begin
				q			<=			16'h0004;
		end
		32'h0000268C: begin
				q			<=			16'h0513;
		end
		32'h0000268E: begin
				q			<=			16'h0010;
		end
		32'h00002690: begin
				q			<=			16'h006F;
		end
		32'h00002692: begin
				q			<=			16'h00C0;
		end
		32'h00002694: begin
				q			<=			16'h00A3;
		end
		32'h00002696: begin
				q			<=			16'h0004;
		end
		32'h00002698: begin
				q			<=			16'h0513;
		end
		32'h0000269A: begin
				q			<=			16'h0010;
		end
		32'h0000269C: begin
				q			<=			16'h2083;
		end
		32'h0000269E: begin
				q			<=			16'h01C1;
		end
		32'h000026A0: begin
				q			<=			16'h2403;
		end
		32'h000026A2: begin
				q			<=			16'h0181;
		end
		32'h000026A4: begin
				q			<=			16'h2483;
		end
		32'h000026A6: begin
				q			<=			16'h0141;
		end
		32'h000026A8: begin
				q			<=			16'h2903;
		end
		32'h000026AA: begin
				q			<=			16'h0101;
		end
		32'h000026AC: begin
				q			<=			16'h2983;
		end
		32'h000026AE: begin
				q			<=			16'h00C1;
		end
		32'h000026B0: begin
				q			<=			16'h2A03;
		end
		32'h000026B2: begin
				q			<=			16'h0081;
		end
		32'h000026B4: begin
				q			<=			16'h2A83;
		end
		32'h000026B6: begin
				q			<=			16'h0041;
		end
		32'h000026B8: begin
				q			<=			16'h2B03;
		end
		32'h000026BA: begin
				q			<=			16'h0001;
		end
		32'h000026BC: begin
				q			<=			16'h0113;
		end
		32'h000026BE: begin
				q			<=			16'h0201;
		end
		32'h000026C0: begin
				q			<=			16'h8067;
		end
		32'h000026C2: begin
				q			<=			16'h0000;
		end
		32'h000026C4: begin
				q			<=			16'h0513;
		end
		32'h000026C6: begin
				q			<=			16'h0000;
		end
		32'h000026C8: begin
				q			<=			16'hF06F;
		end
		32'h000026CA: begin
				q			<=			16'hFD5F;
		end
		32'h000026CC: begin
				q			<=			16'h0513;
		end
		32'h000026CE: begin
				q			<=			16'h0050;
		end
		32'h000026D0: begin
				q			<=			16'hF06F;
		end
		32'h000026D2: begin
				q			<=			16'hFCDF;
		end
		32'h000026D4: begin
				q			<=			16'h0513;
		end
		32'h000026D6: begin
				q			<=			16'h0000;
		end
		32'h000026D8: begin
				q			<=			16'hF06F;
		end
		32'h000026DA: begin
				q			<=			16'hFC5F;
		end
		32'h000026DC: begin
				q			<=			16'h0000;
		end
		32'h000026DE: begin
				q			<=			16'h0000;
		end
		32'h000026E0: begin
				q			<=			16'h17B7;
		end
		32'h000026E2: begin
				q			<=			16'h0001;
		end
		32'h000026E4: begin
				q			<=			16'hA783;
		end
		32'h000026E6: begin
				q			<=			16'hF9C7;
		end
		32'h000026E8: begin
				q			<=			16'h8463;
		end
		32'h000026EA: begin
				q			<=			16'h0607;
		end
		32'h000026EC: begin
				q			<=			16'h0113;
		end
		32'h000026EE: begin
				q			<=			16'hFC01;
		end
		32'h000026F0: begin
				q			<=			16'h2E23;
		end
		32'h000026F2: begin
				q			<=			16'h0211;
		end
		32'h000026F4: begin
				q			<=			16'h2C23;
		end
		32'h000026F6: begin
				q			<=			16'h0281;
		end
		32'h000026F8: begin
				q			<=			16'h8613;
		end
		32'h000026FA: begin
				q			<=			16'h0005;
		end
		32'h000026FC: begin
				q			<=			16'h0413;
		end
		32'h000026FE: begin
				q			<=			16'h0005;
		end
		32'h00002700: begin
				q			<=			16'h0793;
		end
		32'h00002702: begin
				q			<=			16'h0241;
		end
		32'h00002704: begin
				q			<=			16'h2223;
		end
		32'h00002706: begin
				q			<=			16'h00F5;
		end
		32'h00002708: begin
				q			<=			16'h0593;
		end
		32'h0000270A: begin
				q			<=			16'h0041;
		end
		32'h0000270C: begin
				q			<=			16'hF0EF;
		end
		32'h0000270E: begin
				q			<=			16'h9A1F;
		end
		32'h00002710: begin
				q			<=			16'h1863;
		end
		32'h00002712: begin
				q			<=			16'h0205;
		end
		32'h00002714: begin
				q			<=			16'h4783;
		end
		32'h00002716: begin
				q			<=			16'h0041;
		end
		32'h00002718: begin
				q			<=			16'h8063;
		end
		32'h0000271A: begin
				q			<=			16'h0207;
		end
		32'h0000271C: begin
				q			<=			16'h4783;
		end
		32'h0000271E: begin
				q			<=			16'h00F1;
		end
		32'h00002720: begin
				q			<=			16'hF793;
		end
		32'h00002722: begin
				q			<=			16'h0107;
		end
		32'h00002724: begin
				q			<=			16'h0513;
		end
		32'h00002726: begin
				q			<=			16'h0030;
		end
		32'h00002728: begin
				q			<=			16'h8C63;
		end
		32'h0000272A: begin
				q			<=			16'h0007;
		end
		32'h0000272C: begin
				q			<=			16'h0513;
		end
		32'h0000272E: begin
				q			<=			16'h0041;
		end
		32'h00002730: begin
				q			<=			16'hF0EF;
		end
		32'h00002732: begin
				q			<=			16'h931F;
		end
		32'h00002734: begin
				q			<=			16'h2423;
		end
		32'h00002736: begin
				q			<=			16'h00A4;
		end
		32'h00002738: begin
				q			<=			16'h0513;
		end
		32'h0000273A: begin
				q			<=			16'h0004;
		end
		32'h0000273C: begin
				q			<=			16'hF0EF;
		end
		32'h0000273E: begin
				q			<=			16'hDF4F;
		end
		32'h00002740: begin
				q			<=			16'h2083;
		end
		32'h00002742: begin
				q			<=			16'h03C1;
		end
		32'h00002744: begin
				q			<=			16'h2403;
		end
		32'h00002746: begin
				q			<=			16'h0381;
		end
		32'h00002748: begin
				q			<=			16'h0113;
		end
		32'h0000274A: begin
				q			<=			16'h0401;
		end
		32'h0000274C: begin
				q			<=			16'h8067;
		end
		32'h0000274E: begin
				q			<=			16'h0000;
		end
		32'h00002750: begin
				q			<=			16'h0513;
		end
		32'h00002752: begin
				q			<=			16'h0050;
		end
		32'h00002754: begin
				q			<=			16'h8067;
		end
		32'h00002756: begin
				q			<=			16'h0000;
		end
		32'h00002758: begin
				q			<=			16'h0000;
		end
		32'h0000275A: begin
				q			<=			16'h0000;
		end
		32'h0000275C: begin
				q			<=			16'h17B7;
		end
		32'h0000275E: begin
				q			<=			16'h0001;
		end
		32'h00002760: begin
				q			<=			16'hA783;
		end
		32'h00002762: begin
				q			<=			16'hF9C7;
		end
		32'h00002764: begin
				q			<=			16'h8A63;
		end
		32'h00002766: begin
				q			<=			16'h1C07;
		end
		32'h00002768: begin
				q			<=			16'h0113;
		end
		32'h0000276A: begin
				q			<=			16'hFB01;
		end
		32'h0000276C: begin
				q			<=			16'h2623;
		end
		32'h0000276E: begin
				q			<=			16'h0411;
		end
		32'h00002770: begin
				q			<=			16'h2423;
		end
		32'h00002772: begin
				q			<=			16'h0481;
		end
		32'h00002774: begin
				q			<=			16'h2223;
		end
		32'h00002776: begin
				q			<=			16'h0491;
		end
		32'h00002778: begin
				q			<=			16'h2023;
		end
		32'h0000277A: begin
				q			<=			16'h0521;
		end
		32'h0000277C: begin
				q			<=			16'h2E23;
		end
		32'h0000277E: begin
				q			<=			16'h0331;
		end
		32'h00002780: begin
				q			<=			16'h8913;
		end
		32'h00002782: begin
				q			<=			16'h0005;
		end
		32'h00002784: begin
				q			<=			16'h0413;
		end
		32'h00002786: begin
				q			<=			16'h0005;
		end
		32'h00002788: begin
				q			<=			16'h0793;
		end
		32'h0000278A: begin
				q			<=			16'h0241;
		end
		32'h0000278C: begin
				q			<=			16'h2223;
		end
		32'h0000278E: begin
				q			<=			16'h00F5;
		end
		32'h00002790: begin
				q			<=			16'h0513;
		end
		32'h00002792: begin
				q			<=			16'h0030;
		end
		32'h00002794: begin
				q			<=			16'h8863;
		end
		32'h00002796: begin
				q			<=			16'h0005;
		end
		32'h00002798: begin
				q			<=			16'h0493;
		end
		32'h0000279A: begin
				q			<=			16'h0E50;
		end
		32'h0000279C: begin
				q			<=			16'h0993;
		end
		32'h0000279E: begin
				q			<=			16'h02E0;
		end
		32'h000027A0: begin
				q			<=			16'h006F;
		end
		32'h000027A2: begin
				q			<=			16'h01C0;
		end
		32'h000027A4: begin
				q			<=			16'h0513;
		end
		32'h000027A6: begin
				q			<=			16'h0004;
		end
		32'h000027A8: begin
				q			<=			16'hF0EF;
		end
		32'h000027AA: begin
				q			<=			16'hD88F;
		end
		32'h000027AC: begin
				q			<=			16'h006F;
		end
		32'h000027AE: begin
				q			<=			16'h1600;
		end
		32'h000027B0: begin
				q			<=			16'h0513;
		end
		32'h000027B2: begin
				q			<=			16'h0004;
		end
		32'h000027B4: begin
				q			<=			16'hF0EF;
		end
		32'h000027B6: begin
				q			<=			16'hEE4F;
		end
		32'h000027B8: begin
				q			<=			16'h1E63;
		end
		32'h000027BA: begin
				q			<=			16'h0605;
		end
		32'h000027BC: begin
				q			<=			16'h2583;
		end
		32'h000027BE: begin
				q			<=			16'h0104;
		end
		32'h000027C0: begin
				q			<=			16'h8063;
		end
		32'h000027C2: begin
				q			<=			16'h1805;
		end
		32'h000027C4: begin
				q			<=			16'h5603;
		end
		32'h000027C6: begin
				q			<=			16'h0004;
		end
		32'h000027C8: begin
				q			<=			16'h7613;
		end
		32'h000027CA: begin
				q			<=			16'h00F6;
		end
		32'h000027CC: begin
				q			<=			16'h0693;
		end
		32'h000027CE: begin
				q			<=			16'h0200;
		end
		32'h000027D0: begin
				q			<=			16'h1613;
		end
		32'h000027D2: begin
				q			<=			16'h0056;
		end
		32'h000027D4: begin
				q			<=			16'h0513;
		end
		32'h000027D6: begin
				q			<=			16'h0041;
		end
		32'h000027D8: begin
				q			<=			16'hF0EF;
		end
		32'h000027DA: begin
				q			<=			16'hC4CF;
		end
		32'h000027DC: begin
				q			<=			16'h1A63;
		end
		32'h000027DE: begin
				q			<=			16'h0405;
		end
		32'h000027E0: begin
				q			<=			16'h4783;
		end
		32'h000027E2: begin
				q			<=			16'h0041;
		end
		32'h000027E4: begin
				q			<=			16'h8463;
		end
		32'h000027E6: begin
				q			<=			16'h1607;
		end
		32'h000027E8: begin
				q			<=			16'h84E3;
		end
		32'h000027EA: begin
				q			<=			16'hFC97;
		end
		32'h000027EC: begin
				q			<=			16'h82E3;
		end
		32'h000027EE: begin
				q			<=			16'hFD37;
		end
		32'h000027F0: begin
				q			<=			16'h4783;
		end
		32'h000027F2: begin
				q			<=			16'h00F1;
		end
		32'h000027F4: begin
				q			<=			16'hF793;
		end
		32'h000027F6: begin
				q			<=			16'h0087;
		end
		32'h000027F8: begin
				q			<=			16'h9CE3;
		end
		32'h000027FA: begin
				q			<=			16'hFA07;
		end
		32'h000027FC: begin
				q			<=			16'h0713;
		end
		32'h000027FE: begin
				q			<=			16'h0099;
		end
		32'h00002800: begin
				q			<=			16'h2783;
		end
		32'h00002802: begin
				q			<=			16'h0104;
		end
		32'h00002804: begin
				q			<=			16'h0493;
		end
		32'h00002806: begin
				q			<=			16'h0007;
		end
		32'h00002808: begin
				q			<=			16'h8463;
		end
		32'h0000280A: begin
				q			<=			16'h0E07;
		end
		32'h0000280C: begin
				q			<=			16'h4783;
		end
		32'h0000280E: begin
				q			<=			16'h0041;
		end
		32'h00002810: begin
				q			<=			16'h0693;
		end
		32'h00002812: begin
				q			<=			16'h0200;
		end
		32'h00002814: begin
				q			<=			16'h8063;
		end
		32'h00002816: begin
				q			<=			16'h06D7;
		end
		32'h00002818: begin
				q			<=			16'h0693;
		end
		32'h0000281A: begin
				q			<=			16'h0041;
		end
		32'h0000281C: begin
				q			<=			16'h0493;
		end
		32'h0000281E: begin
				q			<=			16'h0119;
		end
		32'h00002820: begin
				q			<=			16'h0613;
		end
		32'h00002822: begin
				q			<=			16'h0050;
		end
		32'h00002824: begin
				q			<=			16'h0513;
		end
		32'h00002826: begin
				q			<=			16'h0E50;
		end
		32'h00002828: begin
				q			<=			16'h0593;
		end
		32'h0000282A: begin
				q			<=			16'h0200;
		end
		32'h0000282C: begin
				q			<=			16'h006F;
		end
		32'h0000282E: begin
				q			<=			16'h0380;
		end
		32'h00002830: begin
				q			<=			16'h0513;
		end
		32'h00002832: begin
				q			<=			16'h0010;
		end
		32'h00002834: begin
				q			<=			16'h2823;
		end
		32'h00002836: begin
				q			<=			16'h0004;
		end
		32'h00002838: begin
				q			<=			16'h0793;
		end
		32'h0000283A: begin
				q			<=			16'h0030;
		end
		32'h0000283C: begin
				q			<=			16'h0A63;
		end
		32'h0000283E: begin
				q			<=			16'h10F5;
		end
		32'h00002840: begin
				q			<=			16'h1663;
		end
		32'h00002842: begin
				q			<=			16'h0C05;
		end
		32'h00002844: begin
				q			<=			16'h0493;
		end
		32'h00002846: begin
				q			<=			16'h0099;
		end
		32'h00002848: begin
				q			<=			16'h006F;
		end
		32'h0000284A: begin
				q			<=			16'h0A80;
		end
		32'h0000284C: begin
				q			<=			16'h0713;
		end
		32'h0000284E: begin
				q			<=			16'h0017;
		end
		32'h00002850: begin
				q			<=			16'h0FA3;
		end
		32'h00002852: begin
				q			<=			16'hFEF7;
		end
		32'h00002854: begin
				q			<=			16'h0063;
		end
		32'h00002856: begin
				q			<=			16'h0297;
		end
		32'h00002858: begin
				q			<=			16'h8693;
		end
		32'h0000285A: begin
				q			<=			16'h0016;
		end
		32'h0000285C: begin
				q			<=			16'hC783;
		end
		32'h0000285E: begin
				q			<=			16'h0006;
		end
		32'h00002860: begin
				q			<=			16'h8863;
		end
		32'h00002862: begin
				q			<=			16'h00B7;
		end
		32'h00002864: begin
				q			<=			16'h94E3;
		end
		32'h00002866: begin
				q			<=			16'hFEC7;
		end
		32'h00002868: begin
				q			<=			16'h0793;
		end
		32'h0000286A: begin
				q			<=			16'h0005;
		end
		32'h0000286C: begin
				q			<=			16'hF06F;
		end
		32'h0000286E: begin
				q			<=			16'hFE1F;
		end
		32'h00002870: begin
				q			<=			16'h0493;
		end
		32'h00002872: begin
				q			<=			16'h0007;
		end
		32'h00002874: begin
				q			<=			16'h4783;
		end
		32'h00002876: begin
				q			<=			16'h00C1;
		end
		32'h00002878: begin
				q			<=			16'h0713;
		end
		32'h0000287A: begin
				q			<=			16'h0200;
		end
		32'h0000287C: begin
				q			<=			16'h8C63;
		end
		32'h0000287E: begin
				q			<=			16'h02E7;
		end
		32'h00002880: begin
				q			<=			16'h0713;
		end
		32'h00002882: begin
				q			<=			16'h02E0;
		end
		32'h00002884: begin
				q			<=			16'h8023;
		end
		32'h00002886: begin
				q			<=			16'h00E4;
		end
		32'h00002888: begin
				q			<=			16'h8693;
		end
		32'h0000288A: begin
				q			<=			16'h0024;
		end
		32'h0000288C: begin
				q			<=			16'h80A3;
		end
		32'h0000288E: begin
				q			<=			16'h00F4;
		end
		32'h00002890: begin
				q			<=			16'h4783;
		end
		32'h00002892: begin
				q			<=			16'h00D1;
		end
		32'h00002894: begin
				q			<=			16'h0713;
		end
		32'h00002896: begin
				q			<=			16'h0200;
		end
		32'h00002898: begin
				q			<=			16'h8863;
		end
		32'h0000289A: begin
				q			<=			16'h08E7;
		end
		32'h0000289C: begin
				q			<=			16'h8693;
		end
		32'h0000289E: begin
				q			<=			16'h0034;
		end
		32'h000028A0: begin
				q			<=			16'h8123;
		end
		32'h000028A2: begin
				q			<=			16'h00F4;
		end
		32'h000028A4: begin
				q			<=			16'h4783;
		end
		32'h000028A6: begin
				q			<=			16'h00E1;
		end
		32'h000028A8: begin
				q			<=			16'h8463;
		end
		32'h000028AA: begin
				q			<=			16'h08E7;
		end
		32'h000028AC: begin
				q			<=			16'h81A3;
		end
		32'h000028AE: begin
				q			<=			16'h00F4;
		end
		32'h000028B0: begin
				q			<=			16'h8493;
		end
		32'h000028B2: begin
				q			<=			16'h0044;
		end
		32'h000028B4: begin
				q			<=			16'h4783;
		end
		32'h000028B6: begin
				q			<=			16'h00F1;
		end
		32'h000028B8: begin
				q			<=			16'h0423;
		end
		32'h000028BA: begin
				q			<=			16'h00F9;
		end
		32'h000028BC: begin
				q			<=			16'h0513;
		end
		32'h000028BE: begin
				q			<=			16'h0201;
		end
		32'h000028C0: begin
				q			<=			16'hF0EF;
		end
		32'h000028C2: begin
				q			<=			16'hC08F;
		end
		32'h000028C4: begin
				q			<=			16'h2023;
		end
		32'h000028C6: begin
				q			<=			16'h00A9;
		end
		32'h000028C8: begin
				q			<=			16'h4783;
		end
		32'h000028CA: begin
				q			<=			16'h01D1;
		end
		32'h000028CC: begin
				q			<=			16'h9793;
		end
		32'h000028CE: begin
				q			<=			16'h0087;
		end
		32'h000028D0: begin
				q			<=			16'h4703;
		end
		32'h000028D2: begin
				q			<=			16'h01C1;
		end
		32'h000028D4: begin
				q			<=			16'hE7B3;
		end
		32'h000028D6: begin
				q			<=			16'h00E7;
		end
		32'h000028D8: begin
				q			<=			16'h1223;
		end
		32'h000028DA: begin
				q			<=			16'h00F9;
		end
		32'h000028DC: begin
				q			<=			16'h4783;
		end
		32'h000028DE: begin
				q			<=			16'h01B1;
		end
		32'h000028E0: begin
				q			<=			16'h9793;
		end
		32'h000028E2: begin
				q			<=			16'h0087;
		end
		32'h000028E4: begin
				q			<=			16'h4703;
		end
		32'h000028E6: begin
				q			<=			16'h01A1;
		end
		32'h000028E8: begin
				q			<=			16'hE7B3;
		end
		32'h000028EA: begin
				q			<=			16'h00E7;
		end
		32'h000028EC: begin
				q			<=			16'h1323;
		end
		32'h000028EE: begin
				q			<=			16'h00F9;
		end
		32'h000028F0: begin
				q			<=			16'h8023;
		end
		32'h000028F2: begin
				q			<=			16'h0004;
		end
		32'h000028F4: begin
				q			<=			16'h0513;
		end
		32'h000028F6: begin
				q			<=			16'h0004;
		end
		32'h000028F8: begin
				q			<=			16'hF0EF;
		end
		32'h000028FA: begin
				q			<=			16'hDA0F;
		end
		32'h000028FC: begin
				q			<=			16'h0793;
		end
		32'h000028FE: begin
				q			<=			16'hFFD5;
		end
		32'h00002900: begin
				q			<=			16'h37B3;
		end
		32'h00002902: begin
				q			<=			16'h00F0;
		end
		32'h00002904: begin
				q			<=			16'h07B3;
		end
		32'h00002906: begin
				q			<=			16'h40F0;
		end
		32'h00002908: begin
				q			<=			16'h7533;
		end
		32'h0000290A: begin
				q			<=			16'h00F5;
		end
		32'h0000290C: begin
				q			<=			16'h2083;
		end
		32'h0000290E: begin
				q			<=			16'h04C1;
		end
		32'h00002910: begin
				q			<=			16'h2403;
		end
		32'h00002912: begin
				q			<=			16'h0481;
		end
		32'h00002914: begin
				q			<=			16'h2483;
		end
		32'h00002916: begin
				q			<=			16'h0441;
		end
		32'h00002918: begin
				q			<=			16'h2903;
		end
		32'h0000291A: begin
				q			<=			16'h0401;
		end
		32'h0000291C: begin
				q			<=			16'h2983;
		end
		32'h0000291E: begin
				q			<=			16'h03C1;
		end
		32'h00002920: begin
				q			<=			16'h0113;
		end
		32'h00002922: begin
				q			<=			16'h0501;
		end
		32'h00002924: begin
				q			<=			16'h8067;
		end
		32'h00002926: begin
				q			<=			16'h0000;
		end
		32'h00002928: begin
				q			<=			16'h8493;
		end
		32'h0000292A: begin
				q			<=			16'h0006;
		end
		32'h0000292C: begin
				q			<=			16'hF06F;
		end
		32'h0000292E: begin
				q			<=			16'hF89F;
		end
		32'h00002930: begin
				q			<=			16'h8493;
		end
		32'h00002932: begin
				q			<=			16'h0006;
		end
		32'h00002934: begin
				q			<=			16'hF06F;
		end
		32'h00002936: begin
				q			<=			16'hF81F;
		end
		32'h00002938: begin
				q			<=			16'h0513;
		end
		32'h0000293A: begin
				q			<=			16'h0050;
		end
		32'h0000293C: begin
				q			<=			16'h8067;
		end
		32'h0000293E: begin
				q			<=			16'h0000;
		end
		32'h00002940: begin
				q			<=			16'h0493;
		end
		32'h00002942: begin
				q			<=			16'h0099;
		end
		32'h00002944: begin
				q			<=			16'h06E3;
		end
		32'h00002946: begin
				q			<=			16'hFA05;
		end
		32'h00002948: begin
				q			<=			16'hF06F;
		end
		32'h0000294A: begin
				q			<=			16'hEEDF;
		end
		32'h0000294C: begin
				q			<=			16'h2823;
		end
		32'h0000294E: begin
				q			<=			16'h0004;
		end
		32'h00002950: begin
				q			<=			16'h0493;
		end
		32'h00002952: begin
				q			<=			16'h0099;
		end
		32'h00002954: begin
				q			<=			16'hF06F;
		end
		32'h00002956: begin
				q			<=			16'hF9DF;
		end
		32'h00002958: begin
				q			<=			16'h0000;
		end
		32'h0000295A: begin
				q			<=			16'h0000;
		end
		32'h0000295C: begin
				q			<=			16'h4063;
		end
		32'h0000295E: begin
				q			<=			16'h0605;
		end
		32'h00002960: begin
				q			<=			16'hC663;
		end
		32'h00002962: begin
				q			<=			16'h0605;
		end
		32'h00002964: begin
				q			<=			16'h8613;
		end
		32'h00002966: begin
				q			<=			16'h0005;
		end
		32'h00002968: begin
				q			<=			16'h0593;
		end
		32'h0000296A: begin
				q			<=			16'h0005;
		end
		32'h0000296C: begin
				q			<=			16'h0513;
		end
		32'h0000296E: begin
				q			<=			16'hFFF0;
		end
		32'h00002970: begin
				q			<=			16'h0C63;
		end
		32'h00002972: begin
				q			<=			16'h0206;
		end
		32'h00002974: begin
				q			<=			16'h0693;
		end
		32'h00002976: begin
				q			<=			16'h0010;
		end
		32'h00002978: begin
				q			<=			16'h7A63;
		end
		32'h0000297A: begin
				q			<=			16'h00B6;
		end
		32'h0000297C: begin
				q			<=			16'h5863;
		end
		32'h0000297E: begin
				q			<=			16'h00C0;
		end
		32'h00002980: begin
				q			<=			16'h1613;
		end
		32'h00002982: begin
				q			<=			16'h0016;
		end
		32'h00002984: begin
				q			<=			16'h9693;
		end
		32'h00002986: begin
				q			<=			16'h0016;
		end
		32'h00002988: begin
				q			<=			16'h6AE3;
		end
		32'h0000298A: begin
				q			<=			16'hFEB6;
		end
		32'h0000298C: begin
				q			<=			16'h0513;
		end
		32'h0000298E: begin
				q			<=			16'h0000;
		end
		32'h00002990: begin
				q			<=			16'hE663;
		end
		32'h00002992: begin
				q			<=			16'h00C5;
		end
		32'h00002994: begin
				q			<=			16'h85B3;
		end
		32'h00002996: begin
				q			<=			16'h40C5;
		end
		32'h00002998: begin
				q			<=			16'h6533;
		end
		32'h0000299A: begin
				q			<=			16'h00D5;
		end
		32'h0000299C: begin
				q			<=			16'hD693;
		end
		32'h0000299E: begin
				q			<=			16'h0016;
		end
		32'h000029A0: begin
				q			<=			16'h5613;
		end
		32'h000029A2: begin
				q			<=			16'h0016;
		end
		32'h000029A4: begin
				q			<=			16'h96E3;
		end
		32'h000029A6: begin
				q			<=			16'hFE06;
		end
		32'h000029A8: begin
				q			<=			16'h8067;
		end
		32'h000029AA: begin
				q			<=			16'h0000;
		end
		32'h000029AC: begin
				q			<=			16'h8293;
		end
		32'h000029AE: begin
				q			<=			16'h0000;
		end
		32'h000029B0: begin
				q			<=			16'hF0EF;
		end
		32'h000029B2: begin
				q			<=			16'hFB5F;
		end
		32'h000029B4: begin
				q			<=			16'h8513;
		end
		32'h000029B6: begin
				q			<=			16'h0005;
		end
		32'h000029B8: begin
				q			<=			16'h8067;
		end
		32'h000029BA: begin
				q			<=			16'h0002;
		end
		32'h000029BC: begin
				q			<=			16'h0533;
		end
		32'h000029BE: begin
				q			<=			16'h40A0;
		end
		32'h000029C0: begin
				q			<=			16'hD863;
		end
		32'h000029C2: begin
				q			<=			16'h0005;
		end
		32'h000029C4: begin
				q			<=			16'h05B3;
		end
		32'h000029C6: begin
				q			<=			16'h40B0;
		end
		32'h000029C8: begin
				q			<=			16'hF06F;
		end
		32'h000029CA: begin
				q			<=			16'hF9DF;
		end
		32'h000029CC: begin
				q			<=			16'h05B3;
		end
		32'h000029CE: begin
				q			<=			16'h40B0;
		end
		32'h000029D0: begin
				q			<=			16'h8293;
		end
		32'h000029D2: begin
				q			<=			16'h0000;
		end
		32'h000029D4: begin
				q			<=			16'hF0EF;
		end
		32'h000029D6: begin
				q			<=			16'hF91F;
		end
		32'h000029D8: begin
				q			<=			16'h0533;
		end
		32'h000029DA: begin
				q			<=			16'h40A0;
		end
		32'h000029DC: begin
				q			<=			16'h8067;
		end
		32'h000029DE: begin
				q			<=			16'h0002;
		end
		32'h000029E0: begin
				q			<=			16'h8293;
		end
		32'h000029E2: begin
				q			<=			16'h0000;
		end
		32'h000029E4: begin
				q			<=			16'hCA63;
		end
		32'h000029E6: begin
				q			<=			16'h0005;
		end
		32'h000029E8: begin
				q			<=			16'h4C63;
		end
		32'h000029EA: begin
				q			<=			16'h0005;
		end
		32'h000029EC: begin
				q			<=			16'hF0EF;
		end
		32'h000029EE: begin
				q			<=			16'hF79F;
		end
		32'h000029F0: begin
				q			<=			16'h8513;
		end
		32'h000029F2: begin
				q			<=			16'h0005;
		end
		32'h000029F4: begin
				q			<=			16'h8067;
		end
		32'h000029F6: begin
				q			<=			16'h0002;
		end
		32'h000029F8: begin
				q			<=			16'h05B3;
		end
		32'h000029FA: begin
				q			<=			16'h40B0;
		end
		32'h000029FC: begin
				q			<=			16'h58E3;
		end
		32'h000029FE: begin
				q			<=			16'hFE05;
		end
		32'h00002A00: begin
				q			<=			16'h0533;
		end
		32'h00002A02: begin
				q			<=			16'h40A0;
		end
		32'h00002A04: begin
				q			<=			16'hF0EF;
		end
		32'h00002A06: begin
				q			<=			16'hF61F;
		end
		32'h00002A08: begin
				q			<=			16'h0533;
		end
		32'h00002A0A: begin
				q			<=			16'h40B0;
		end
		32'h00002A0C: begin
				q			<=			16'h8067;
		end
		32'h00002A0E: begin
				q			<=			16'h0002;
		end
		32'h00002A10: begin
				q			<=			16'h0000;
		end
		32'h00002A12: begin
				q			<=			16'h0000;
		end
		32'h00002A14: begin
				q			<=			16'h0613;
		end
		32'h00002A16: begin
				q			<=			16'h0005;
		end
		32'h00002A18: begin
				q			<=			16'h0513;
		end
		32'h00002A1A: begin
				q			<=			16'h0000;
		end
		32'h00002A1C: begin
				q			<=			16'hF693;
		end
		32'h00002A1E: begin
				q			<=			16'h0015;
		end
		32'h00002A20: begin
				q			<=			16'h8463;
		end
		32'h00002A22: begin
				q			<=			16'h0006;
		end
		32'h00002A24: begin
				q			<=			16'h0533;
		end
		32'h00002A26: begin
				q			<=			16'h00C5;
		end
		32'h00002A28: begin
				q			<=			16'hD593;
		end
		32'h00002A2A: begin
				q			<=			16'h0015;
		end
		32'h00002A2C: begin
				q			<=			16'h1613;
		end
		32'h00002A2E: begin
				q			<=			16'h0016;
		end
		32'h00002A30: begin
				q			<=			16'h96E3;
		end
		32'h00002A32: begin
				q			<=			16'hFE05;
		end
		32'h00002A34: begin
				q			<=			16'h8067;
		end
		32'h00002A36: begin
				q			<=			16'h0000;
		end
		32'h00002A38: begin
				q			<=			16'h0000;
		end
		32'h00002A3A: begin
				q			<=			16'h0000;
		end
		32'h00002A3C: begin
				q			<=			16'h0113;
		end
		32'h00002A3E: begin
				q			<=			16'hFC01;
		end
		32'h00002A40: begin
				q			<=			16'h0313;
		end
		32'h00002A42: begin
				q			<=			16'h0000;
		end
		32'h00002A44: begin
				q			<=			16'h2623;
		end
		32'h00002A46: begin
				q			<=			16'h01B1;
		end
		32'h00002A48: begin
				q			<=			16'h006F;
		end
		32'h00002A4A: begin
				q			<=			16'h00C0;
		end
		32'h00002A4C: begin
				q			<=			16'h0113;
		end
		32'h00002A4E: begin
				q			<=			16'hFC01;
		end
		32'h00002A50: begin
				q			<=			16'h0313;
		end
		32'h00002A52: begin
				q			<=			16'hFF00;
		end
		32'h00002A54: begin
				q			<=			16'h2823;
		end
		32'h00002A56: begin
				q			<=			16'h01A1;
		end
		32'h00002A58: begin
				q			<=			16'h2A23;
		end
		32'h00002A5A: begin
				q			<=			16'h0191;
		end
		32'h00002A5C: begin
				q			<=			16'h2C23;
		end
		32'h00002A5E: begin
				q			<=			16'h0181;
		end
		32'h00002A60: begin
				q			<=			16'h2E23;
		end
		32'h00002A62: begin
				q			<=			16'h0171;
		end
		32'h00002A64: begin
				q			<=			16'h006F;
		end
		32'h00002A66: begin
				q			<=			16'h00C0;
		end
		32'h00002A68: begin
				q			<=			16'h0113;
		end
		32'h00002A6A: begin
				q			<=			16'hFC01;
		end
		32'h00002A6C: begin
				q			<=			16'h0313;
		end
		32'h00002A6E: begin
				q			<=			16'hFE00;
		end
		32'h00002A70: begin
				q			<=			16'h2023;
		end
		32'h00002A72: begin
				q			<=			16'h0361;
		end
		32'h00002A74: begin
				q			<=			16'h2223;
		end
		32'h00002A76: begin
				q			<=			16'h0351;
		end
		32'h00002A78: begin
				q			<=			16'h2423;
		end
		32'h00002A7A: begin
				q			<=			16'h0341;
		end
		32'h00002A7C: begin
				q			<=			16'h2623;
		end
		32'h00002A7E: begin
				q			<=			16'h0331;
		end
		32'h00002A80: begin
				q			<=			16'h2823;
		end
		32'h00002A82: begin
				q			<=			16'h0321;
		end
		32'h00002A84: begin
				q			<=			16'h2A23;
		end
		32'h00002A86: begin
				q			<=			16'h0291;
		end
		32'h00002A88: begin
				q			<=			16'h2C23;
		end
		32'h00002A8A: begin
				q			<=			16'h0281;
		end
		32'h00002A8C: begin
				q			<=			16'h2E23;
		end
		32'h00002A8E: begin
				q			<=			16'h0211;
		end
		32'h00002A90: begin
				q			<=			16'h0133;
		end
		32'h00002A92: begin
				q			<=			16'h4061;
		end
		32'h00002A94: begin
				q			<=			16'h8067;
		end
		32'h00002A96: begin
				q			<=			16'h0002;
		end
		32'h00002A98: begin
				q			<=			16'h0113;
		end
		32'h00002A9A: begin
				q			<=			16'hFF01;
		end
		32'h00002A9C: begin
				q			<=			16'h2023;
		end
		32'h00002A9E: begin
				q			<=			16'h0121;
		end
		32'h00002AA0: begin
				q			<=			16'h2223;
		end
		32'h00002AA2: begin
				q			<=			16'h0091;
		end
		32'h00002AA4: begin
				q			<=			16'h2423;
		end
		32'h00002AA6: begin
				q			<=			16'h0081;
		end
		32'h00002AA8: begin
				q			<=			16'h2623;
		end
		32'h00002AAA: begin
				q			<=			16'h0011;
		end
		32'h00002AAC: begin
				q			<=			16'h8067;
		end
		32'h00002AAE: begin
				q			<=			16'h0002;
		end
		32'h00002AB0: begin
				q			<=			16'h2D83;
		end
		32'h00002AB2: begin
				q			<=			16'h00C1;
		end
		32'h00002AB4: begin
				q			<=			16'h0113;
		end
		32'h00002AB6: begin
				q			<=			16'h0101;
		end
		32'h00002AB8: begin
				q			<=			16'h2D03;
		end
		32'h00002ABA: begin
				q			<=			16'h0001;
		end
		32'h00002ABC: begin
				q			<=			16'h2C83;
		end
		32'h00002ABE: begin
				q			<=			16'h0041;
		end
		32'h00002AC0: begin
				q			<=			16'h2C03;
		end
		32'h00002AC2: begin
				q			<=			16'h0081;
		end
		32'h00002AC4: begin
				q			<=			16'h2B83;
		end
		32'h00002AC6: begin
				q			<=			16'h00C1;
		end
		32'h00002AC8: begin
				q			<=			16'h0113;
		end
		32'h00002ACA: begin
				q			<=			16'h0101;
		end
		32'h00002ACC: begin
				q			<=			16'h2B03;
		end
		32'h00002ACE: begin
				q			<=			16'h0001;
		end
		32'h00002AD0: begin
				q			<=			16'h2A83;
		end
		32'h00002AD2: begin
				q			<=			16'h0041;
		end
		32'h00002AD4: begin
				q			<=			16'h2A03;
		end
		32'h00002AD6: begin
				q			<=			16'h0081;
		end
		32'h00002AD8: begin
				q			<=			16'h2983;
		end
		32'h00002ADA: begin
				q			<=			16'h00C1;
		end
		32'h00002ADC: begin
				q			<=			16'h0113;
		end
		32'h00002ADE: begin
				q			<=			16'h0101;
		end
		32'h00002AE0: begin
				q			<=			16'h2903;
		end
		32'h00002AE2: begin
				q			<=			16'h0001;
		end
		32'h00002AE4: begin
				q			<=			16'h2483;
		end
		32'h00002AE6: begin
				q			<=			16'h0041;
		end
		32'h00002AE8: begin
				q			<=			16'h2403;
		end
		32'h00002AEA: begin
				q			<=			16'h0081;
		end
		32'h00002AEC: begin
				q			<=			16'h2083;
		end
		32'h00002AEE: begin
				q			<=			16'h00C1;
		end
		32'h00002AF0: begin
				q			<=			16'h0113;
		end
		32'h00002AF2: begin
				q			<=			16'h0101;
		end
		32'h00002AF4: begin
				q			<=			16'h8067;
		end
		32'h00002AF6: begin
				q			<=			16'h0000;
		end
		32'h00002AF8: begin
				q			<=			16'hC7B3;
		end
		32'h00002AFA: begin
				q			<=			16'h00A5;
		end
		32'h00002AFC: begin
				q			<=			16'hF793;
		end
		32'h00002AFE: begin
				q			<=			16'h0037;
		end
		32'h00002B00: begin
				q			<=			16'h0733;
		end
		32'h00002B02: begin
				q			<=			16'h00C5;
		end
		32'h00002B04: begin
				q			<=			16'h9663;
		end
		32'h00002B06: begin
				q			<=			16'h0007;
		end
		32'h00002B08: begin
				q			<=			16'h0793;
		end
		32'h00002B0A: begin
				q			<=			16'h0030;
		end
		32'h00002B0C: begin
				q			<=			16'hE463;
		end
		32'h00002B0E: begin
				q			<=			16'h02C7;
		end
		32'h00002B10: begin
				q			<=			16'h0793;
		end
		32'h00002B12: begin
				q			<=			16'h0005;
		end
		32'h00002B14: begin
				q			<=			16'h6C63;
		end
		32'h00002B16: begin
				q			<=			16'h00E5;
		end
		32'h00002B18: begin
				q			<=			16'h8067;
		end
		32'h00002B1A: begin
				q			<=			16'h0000;
		end
		32'h00002B1C: begin
				q			<=			16'hC683;
		end
		32'h00002B1E: begin
				q			<=			16'h0005;
		end
		32'h00002B20: begin
				q			<=			16'h8793;
		end
		32'h00002B22: begin
				q			<=			16'h0017;
		end
		32'h00002B24: begin
				q			<=			16'h8593;
		end
		32'h00002B26: begin
				q			<=			16'h0015;
		end
		32'h00002B28: begin
				q			<=			16'h8FA3;
		end
		32'h00002B2A: begin
				q			<=			16'hFED7;
		end
		32'h00002B2C: begin
				q			<=			16'hE8E3;
		end
		32'h00002B2E: begin
				q			<=			16'hFEE7;
		end
		32'h00002B30: begin
				q			<=			16'h8067;
		end
		32'h00002B32: begin
				q			<=			16'h0000;
		end
		32'h00002B34: begin
				q			<=			16'h7793;
		end
		32'h00002B36: begin
				q			<=			16'h0035;
		end
		32'h00002B38: begin
				q			<=			16'h9263;
		end
		32'h00002B3A: begin
				q			<=			16'h0807;
		end
		32'h00002B3C: begin
				q			<=			16'h0793;
		end
		32'h00002B3E: begin
				q			<=			16'h0005;
		end
		32'h00002B40: begin
				q			<=			16'h7693;
		end
		32'h00002B42: begin
				q			<=			16'hFFC7;
		end
		32'h00002B44: begin
				q			<=			16'h8613;
		end
		32'h00002B46: begin
				q			<=			16'hFE06;
		end
		32'h00002B48: begin
				q			<=			16'hF663;
		end
		32'h00002B4A: begin
				q			<=			16'h08C7;
		end
		32'h00002B4C: begin
				q			<=			16'hA383;
		end
		32'h00002B4E: begin
				q			<=			16'h0005;
		end
		32'h00002B50: begin
				q			<=			16'hA283;
		end
		32'h00002B52: begin
				q			<=			16'h0045;
		end
		32'h00002B54: begin
				q			<=			16'hAF83;
		end
		32'h00002B56: begin
				q			<=			16'h0085;
		end
		32'h00002B58: begin
				q			<=			16'hAF03;
		end
		32'h00002B5A: begin
				q			<=			16'h00C5;
		end
		32'h00002B5C: begin
				q			<=			16'hAE83;
		end
		32'h00002B5E: begin
				q			<=			16'h0105;
		end
		32'h00002B60: begin
				q			<=			16'hAE03;
		end
		32'h00002B62: begin
				q			<=			16'h0145;
		end
		32'h00002B64: begin
				q			<=			16'hA303;
		end
		32'h00002B66: begin
				q			<=			16'h0185;
		end
		32'h00002B68: begin
				q			<=			16'hA883;
		end
		32'h00002B6A: begin
				q			<=			16'h01C5;
		end
		32'h00002B6C: begin
				q			<=			16'h8593;
		end
		32'h00002B6E: begin
				q			<=			16'h0245;
		end
		32'h00002B70: begin
				q			<=			16'h8793;
		end
		32'h00002B72: begin
				q			<=			16'h0247;
		end
		32'h00002B74: begin
				q			<=			16'hA803;
		end
		32'h00002B76: begin
				q			<=			16'hFFC5;
		end
		32'h00002B78: begin
				q			<=			16'hAE23;
		end
		32'h00002B7A: begin
				q			<=			16'hFC77;
		end
		32'h00002B7C: begin
				q			<=			16'hA023;
		end
		32'h00002B7E: begin
				q			<=			16'hFE57;
		end
		32'h00002B80: begin
				q			<=			16'hA223;
		end
		32'h00002B82: begin
				q			<=			16'hFFF7;
		end
		32'h00002B84: begin
				q			<=			16'hA423;
		end
		32'h00002B86: begin
				q			<=			16'hFFE7;
		end
		32'h00002B88: begin
				q			<=			16'hA623;
		end
		32'h00002B8A: begin
				q			<=			16'hFFD7;
		end
		32'h00002B8C: begin
				q			<=			16'hA823;
		end
		32'h00002B8E: begin
				q			<=			16'hFFC7;
		end
		32'h00002B90: begin
				q			<=			16'hAA23;
		end
		32'h00002B92: begin
				q			<=			16'hFE67;
		end
		32'h00002B94: begin
				q			<=			16'hAC23;
		end
		32'h00002B96: begin
				q			<=			16'hFF17;
		end
		32'h00002B98: begin
				q			<=			16'hAE23;
		end
		32'h00002B9A: begin
				q			<=			16'hFF07;
		end
		32'h00002B9C: begin
				q			<=			16'hF06F;
		end
		32'h00002B9E: begin
				q			<=			16'hFADF;
		end
		32'h00002BA0: begin
				q			<=			16'hC683;
		end
		32'h00002BA2: begin
				q			<=			16'h0005;
		end
		32'h00002BA4: begin
				q			<=			16'h8793;
		end
		32'h00002BA6: begin
				q			<=			16'h0017;
		end
		32'h00002BA8: begin
				q			<=			16'h8593;
		end
		32'h00002BAA: begin
				q			<=			16'h0015;
		end
		32'h00002BAC: begin
				q			<=			16'h8FA3;
		end
		32'h00002BAE: begin
				q			<=			16'hFED7;
		end
		32'h00002BB0: begin
				q			<=			16'hF693;
		end
		32'h00002BB2: begin
				q			<=			16'h0037;
		end
		32'h00002BB4: begin
				q			<=			16'h96E3;
		end
		32'h00002BB6: begin
				q			<=			16'hFE06;
		end
		32'h00002BB8: begin
				q			<=			16'hF06F;
		end
		32'h00002BBA: begin
				q			<=			16'hF89F;
		end
		32'h00002BBC: begin
				q			<=			16'h0793;
		end
		32'h00002BBE: begin
				q			<=			16'h0005;
		end
		32'h00002BC0: begin
				q			<=			16'hF06F;
		end
		32'h00002BC2: begin
				q			<=			16'hFF1F;
		end
		32'h00002BC4: begin
				q			<=			16'hA603;
		end
		32'h00002BC6: begin
				q			<=			16'h0005;
		end
		32'h00002BC8: begin
				q			<=			16'h8793;
		end
		32'h00002BCA: begin
				q			<=			16'h0047;
		end
		32'h00002BCC: begin
				q			<=			16'h8593;
		end
		32'h00002BCE: begin
				q			<=			16'h0045;
		end
		32'h00002BD0: begin
				q			<=			16'hAE23;
		end
		32'h00002BD2: begin
				q			<=			16'hFEC7;
		end
		32'h00002BD4: begin
				q			<=			16'hE8E3;
		end
		32'h00002BD6: begin
				q			<=			16'hFED7;
		end
		32'h00002BD8: begin
				q			<=			16'hEAE3;
		end
		32'h00002BDA: begin
				q			<=			16'hF4E7;
		end
		32'h00002BDC: begin
				q			<=			16'h8067;
		end
		32'h00002BDE: begin
				q			<=			16'h0000;
		end
		32'h00002BE0: begin
				q			<=			16'h0000;
		end
		32'h00002BE2: begin
				q			<=			16'h0000;
		end
		32'h00002BE4: begin
				q			<=			16'h0813;
		end
		32'h00002BE6: begin
				q			<=			16'h00F0;
		end
		32'h00002BE8: begin
				q			<=			16'h0713;
		end
		32'h00002BEA: begin
				q			<=			16'h0005;
		end
		32'h00002BEC: begin
				q			<=			16'h7E63;
		end
		32'h00002BEE: begin
				q			<=			16'h02C8;
		end
		32'h00002BF0: begin
				q			<=			16'h7793;
		end
		32'h00002BF2: begin
				q			<=			16'h00F7;
		end
		32'h00002BF4: begin
				q			<=			16'h9063;
		end
		32'h00002BF6: begin
				q			<=			16'h0A07;
		end
		32'h00002BF8: begin
				q			<=			16'h9263;
		end
		32'h00002BFA: begin
				q			<=			16'h0805;
		end
		32'h00002BFC: begin
				q			<=			16'h7693;
		end
		32'h00002BFE: begin
				q			<=			16'hFF06;
		end
		32'h00002C00: begin
				q			<=			16'h7613;
		end
		32'h00002C02: begin
				q			<=			16'h00F6;
		end
		32'h00002C04: begin
				q			<=			16'h86B3;
		end
		32'h00002C06: begin
				q			<=			16'h00E6;
		end
		32'h00002C08: begin
				q			<=			16'h2023;
		end
		32'h00002C0A: begin
				q			<=			16'h00B7;
		end
		32'h00002C0C: begin
				q			<=			16'h2223;
		end
		32'h00002C0E: begin
				q			<=			16'h00B7;
		end
		32'h00002C10: begin
				q			<=			16'h2423;
		end
		32'h00002C12: begin
				q			<=			16'h00B7;
		end
		32'h00002C14: begin
				q			<=			16'h2623;
		end
		32'h00002C16: begin
				q			<=			16'h00B7;
		end
		32'h00002C18: begin
				q			<=			16'h0713;
		end
		32'h00002C1A: begin
				q			<=			16'h0107;
		end
		32'h00002C1C: begin
				q			<=			16'h66E3;
		end
		32'h00002C1E: begin
				q			<=			16'hFED7;
		end
		32'h00002C20: begin
				q			<=			16'h1463;
		end
		32'h00002C22: begin
				q			<=			16'h0006;
		end
		32'h00002C24: begin
				q			<=			16'h8067;
		end
		32'h00002C26: begin
				q			<=			16'h0000;
		end
		32'h00002C28: begin
				q			<=			16'h06B3;
		end
		32'h00002C2A: begin
				q			<=			16'h40C8;
		end
		32'h00002C2C: begin
				q			<=			16'h9693;
		end
		32'h00002C2E: begin
				q			<=			16'h0026;
		end
		32'h00002C30: begin
				q			<=			16'h0297;
		end
		32'h00002C32: begin
				q			<=			16'h0000;
		end
		32'h00002C34: begin
				q			<=			16'h86B3;
		end
		32'h00002C36: begin
				q			<=			16'h0056;
		end
		32'h00002C38: begin
				q			<=			16'h8067;
		end
		32'h00002C3A: begin
				q			<=			16'h00C6;
		end
		32'h00002C3C: begin
				q			<=			16'h0723;
		end
		32'h00002C3E: begin
				q			<=			16'h00B7;
		end
		32'h00002C40: begin
				q			<=			16'h06A3;
		end
		32'h00002C42: begin
				q			<=			16'h00B7;
		end
		32'h00002C44: begin
				q			<=			16'h0623;
		end
		32'h00002C46: begin
				q			<=			16'h00B7;
		end
		32'h00002C48: begin
				q			<=			16'h05A3;
		end
		32'h00002C4A: begin
				q			<=			16'h00B7;
		end
		32'h00002C4C: begin
				q			<=			16'h0523;
		end
		32'h00002C4E: begin
				q			<=			16'h00B7;
		end
		32'h00002C50: begin
				q			<=			16'h04A3;
		end
		32'h00002C52: begin
				q			<=			16'h00B7;
		end
		32'h00002C54: begin
				q			<=			16'h0423;
		end
		32'h00002C56: begin
				q			<=			16'h00B7;
		end
		32'h00002C58: begin
				q			<=			16'h03A3;
		end
		32'h00002C5A: begin
				q			<=			16'h00B7;
		end
		32'h00002C5C: begin
				q			<=			16'h0323;
		end
		32'h00002C5E: begin
				q			<=			16'h00B7;
		end
		32'h00002C60: begin
				q			<=			16'h02A3;
		end
		32'h00002C62: begin
				q			<=			16'h00B7;
		end
		32'h00002C64: begin
				q			<=			16'h0223;
		end
		32'h00002C66: begin
				q			<=			16'h00B7;
		end
		32'h00002C68: begin
				q			<=			16'h01A3;
		end
		32'h00002C6A: begin
				q			<=			16'h00B7;
		end
		32'h00002C6C: begin
				q			<=			16'h0123;
		end
		32'h00002C6E: begin
				q			<=			16'h00B7;
		end
		32'h00002C70: begin
				q			<=			16'h00A3;
		end
		32'h00002C72: begin
				q			<=			16'h00B7;
		end
		32'h00002C74: begin
				q			<=			16'h0023;
		end
		32'h00002C76: begin
				q			<=			16'h00B7;
		end
		32'h00002C78: begin
				q			<=			16'h8067;
		end
		32'h00002C7A: begin
				q			<=			16'h0000;
		end
		32'h00002C7C: begin
				q			<=			16'hF593;
		end
		32'h00002C7E: begin
				q			<=			16'h0FF5;
		end
		32'h00002C80: begin
				q			<=			16'h9693;
		end
		32'h00002C82: begin
				q			<=			16'h0085;
		end
		32'h00002C84: begin
				q			<=			16'hE5B3;
		end
		32'h00002C86: begin
				q			<=			16'h00D5;
		end
		32'h00002C88: begin
				q			<=			16'h9693;
		end
		32'h00002C8A: begin
				q			<=			16'h0105;
		end
		32'h00002C8C: begin
				q			<=			16'hE5B3;
		end
		32'h00002C8E: begin
				q			<=			16'h00D5;
		end
		32'h00002C90: begin
				q			<=			16'hF06F;
		end
		32'h00002C92: begin
				q			<=			16'hF6DF;
		end
		32'h00002C94: begin
				q			<=			16'h9693;
		end
		32'h00002C96: begin
				q			<=			16'h0027;
		end
		32'h00002C98: begin
				q			<=			16'h0297;
		end
		32'h00002C9A: begin
				q			<=			16'h0000;
		end
		32'h00002C9C: begin
				q			<=			16'h86B3;
		end
		32'h00002C9E: begin
				q			<=			16'h0056;
		end
		32'h00002CA0: begin
				q			<=			16'h8293;
		end
		32'h00002CA2: begin
				q			<=			16'h0000;
		end
		32'h00002CA4: begin
				q			<=			16'h80E7;
		end
		32'h00002CA6: begin
				q			<=			16'hFA06;
		end
		32'h00002CA8: begin
				q			<=			16'h8093;
		end
		32'h00002CAA: begin
				q			<=			16'h0002;
		end
		32'h00002CAC: begin
				q			<=			16'h8793;
		end
		32'h00002CAE: begin
				q			<=			16'hFF07;
		end
		32'h00002CB0: begin
				q			<=			16'h0733;
		end
		32'h00002CB2: begin
				q			<=			16'h40F7;
		end
		32'h00002CB4: begin
				q			<=			16'h0633;
		end
		32'h00002CB6: begin
				q			<=			16'h00F6;
		end
		32'h00002CB8: begin
				q			<=			16'h78E3;
		end
		32'h00002CBA: begin
				q			<=			16'hF6C8;
		end
		32'h00002CBC: begin
				q			<=			16'hF06F;
		end
		32'h00002CBE: begin
				q			<=			16'hF3DF;
		end
		32'h00002CC0: begin
				q			<=			16'h0113;
		end
		32'h00002CC2: begin
				q			<=			16'hF701;
		end
		32'h00002CC4: begin
				q			<=			16'h2E23;
		end
		32'h00002CC6: begin
				q			<=			16'h0611;
		end
		32'h00002CC8: begin
				q			<=			16'h2C23;
		end
		32'h00002CCA: begin
				q			<=			16'h0681;
		end
		32'h00002CCC: begin
				q			<=			16'h2A23;
		end
		32'h00002CCE: begin
				q			<=			16'h0691;
		end
		32'h00002CD0: begin
				q			<=			16'h2023;
		end
		32'h00002CD2: begin
				q			<=			16'h08E1;
		end
		32'h00002CD4: begin
				q			<=			16'h2223;
		end
		32'h00002CD6: begin
				q			<=			16'h08F1;
		end
		32'h00002CD8: begin
				q			<=			16'h2423;
		end
		32'h00002CDA: begin
				q			<=			16'h0901;
		end
		32'h00002CDC: begin
				q			<=			16'h2623;
		end
		32'h00002CDE: begin
				q			<=			16'h0911;
		end
		32'h00002CE0: begin
				q			<=			16'h5263;
		end
		32'h00002CE2: begin
				q			<=			16'h0206;
		end
		32'h00002CE4: begin
				q			<=			16'h0793;
		end
		32'h00002CE6: begin
				q			<=			16'h08B0;
		end
		32'h00002CE8: begin
				q			<=			16'h2023;
		end
		32'h00002CEA: begin
				q			<=			16'h00F5;
		end
		32'h00002CEC: begin
				q			<=			16'h0513;
		end
		32'h00002CEE: begin
				q			<=			16'hFFF0;
		end
		32'h00002CF0: begin
				q			<=			16'h2083;
		end
		32'h00002CF2: begin
				q			<=			16'h07C1;
		end
		32'h00002CF4: begin
				q			<=			16'h2403;
		end
		32'h00002CF6: begin
				q			<=			16'h0781;
		end
		32'h00002CF8: begin
				q			<=			16'h2483;
		end
		32'h00002CFA: begin
				q			<=			16'h0741;
		end
		32'h00002CFC: begin
				q			<=			16'h0113;
		end
		32'h00002CFE: begin
				q			<=			16'h0901;
		end
		32'h00002D00: begin
				q			<=			16'h8067;
		end
		32'h00002D02: begin
				q			<=			16'h0000;
		end
		32'h00002D04: begin
				q			<=			16'h0793;
		end
		32'h00002D06: begin
				q			<=			16'h2080;
		end
		32'h00002D08: begin
				q			<=			16'h1A23;
		end
		32'h00002D0A: begin
				q			<=			16'h00F1;
		end
		32'h00002D0C: begin
				q			<=			16'h2423;
		end
		32'h00002D0E: begin
				q			<=			16'h00B1;
		end
		32'h00002D10: begin
				q			<=			16'h2C23;
		end
		32'h00002D12: begin
				q			<=			16'h00B1;
		end
		32'h00002D14: begin
				q			<=			16'h0413;
		end
		32'h00002D16: begin
				q			<=			16'h0006;
		end
		32'h00002D18: begin
				q			<=			16'h0793;
		end
		32'h00002D1A: begin
				q			<=			16'h0000;
		end
		32'h00002D1C: begin
				q			<=			16'h0463;
		end
		32'h00002D1E: begin
				q			<=			16'h0006;
		end
		32'h00002D20: begin
				q			<=			16'h0793;
		end
		32'h00002D22: begin
				q			<=			16'hFFF6;
		end
		32'h00002D24: begin
				q			<=			16'h8613;
		end
		32'h00002D26: begin
				q			<=			16'h0006;
		end
		32'h00002D28: begin
				q			<=			16'h2823;
		end
		32'h00002D2A: begin
				q			<=			16'h00F1;
		end
		32'h00002D2C: begin
				q			<=			16'h2E23;
		end
		32'h00002D2E: begin
				q			<=			16'h00F1;
		end
		32'h00002D30: begin
				q			<=			16'h0693;
		end
		32'h00002D32: begin
				q			<=			16'h0801;
		end
		32'h00002D34: begin
				q			<=			16'h0793;
		end
		32'h00002D36: begin
				q			<=			16'hFFF0;
		end
		32'h00002D38: begin
				q			<=			16'h0593;
		end
		32'h00002D3A: begin
				q			<=			16'h0081;
		end
		32'h00002D3C: begin
				q			<=			16'h1B23;
		end
		32'h00002D3E: begin
				q			<=			16'h00F1;
		end
		32'h00002D40: begin
				q			<=			16'h0493;
		end
		32'h00002D42: begin
				q			<=			16'h0005;
		end
		32'h00002D44: begin
				q			<=			16'h2223;
		end
		32'h00002D46: begin
				q			<=			16'h00D1;
		end
		32'h00002D48: begin
				q			<=			16'h00EF;
		end
		32'h00002D4A: begin
				q			<=			16'h1900;
		end
		32'h00002D4C: begin
				q			<=			16'h0793;
		end
		32'h00002D4E: begin
				q			<=			16'hFFF0;
		end
		32'h00002D50: begin
				q			<=			16'h5663;
		end
		32'h00002D52: begin
				q			<=			16'h00F5;
		end
		32'h00002D54: begin
				q			<=			16'h0793;
		end
		32'h00002D56: begin
				q			<=			16'h08B0;
		end
		32'h00002D58: begin
				q			<=			16'hA023;
		end
		32'h00002D5A: begin
				q			<=			16'h00F4;
		end
		32'h00002D5C: begin
				q			<=			16'h0AE3;
		end
		32'h00002D5E: begin
				q			<=			16'hF804;
		end
		32'h00002D60: begin
				q			<=			16'h2783;
		end
		32'h00002D62: begin
				q			<=			16'h0081;
		end
		32'h00002D64: begin
				q			<=			16'h8023;
		end
		32'h00002D66: begin
				q			<=			16'h0007;
		end
		32'h00002D68: begin
				q			<=			16'hF06F;
		end
		32'h00002D6A: begin
				q			<=			16'hF89F;
		end
		32'h00002D6C: begin
				q			<=			16'h0113;
		end
		32'h00002D6E: begin
				q			<=			16'hF601;
		end
		32'h00002D70: begin
				q			<=			16'h2A23;
		end
		32'h00002D72: begin
				q			<=			16'h08F1;
		end
		32'h00002D74: begin
				q			<=			16'h2A23;
		end
		32'h00002D76: begin
				q			<=			16'h0691;
		end
		32'h00002D78: begin
				q			<=			16'h2623;
		end
		32'h00002D7A: begin
				q			<=			16'h08D1;
		end
		32'h00002D7C: begin
				q			<=			16'h2823;
		end
		32'h00002D7E: begin
				q			<=			16'h08E1;
		end
		32'h00002D80: begin
				q			<=			16'h2C23;
		end
		32'h00002D82: begin
				q			<=			16'h0901;
		end
		32'h00002D84: begin
				q			<=			16'h2E23;
		end
		32'h00002D86: begin
				q			<=			16'h0911;
		end
		32'h00002D88: begin
				q			<=			16'hE797;
		end
		32'h00002D8A: begin
				q			<=			16'h0000;
		end
		32'h00002D8C: begin
				q			<=			16'h8793;
		end
		32'h00002D8E: begin
				q			<=			16'hB507;
		end
		32'h00002D90: begin
				q			<=			16'h2E23;
		end
		32'h00002D92: begin
				q			<=			16'h0611;
		end
		32'h00002D94: begin
				q			<=			16'h2C23;
		end
		32'h00002D96: begin
				q			<=			16'h0681;
		end
		32'h00002D98: begin
				q			<=			16'hA483;
		end
		32'h00002D9A: begin
				q			<=			16'h0007;
		end
		32'h00002D9C: begin
				q			<=			16'hD263;
		end
		32'h00002D9E: begin
				q			<=			16'h0205;
		end
		32'h00002DA0: begin
				q			<=			16'h0793;
		end
		32'h00002DA2: begin
				q			<=			16'h08B0;
		end
		32'h00002DA4: begin
				q			<=			16'hA023;
		end
		32'h00002DA6: begin
				q			<=			16'h00F4;
		end
		32'h00002DA8: begin
				q			<=			16'h0513;
		end
		32'h00002DAA: begin
				q			<=			16'hFFF0;
		end
		32'h00002DAC: begin
				q			<=			16'h2083;
		end
		32'h00002DAE: begin
				q			<=			16'h07C1;
		end
		32'h00002DB0: begin
				q			<=			16'h2403;
		end
		32'h00002DB2: begin
				q			<=			16'h0781;
		end
		32'h00002DB4: begin
				q			<=			16'h2483;
		end
		32'h00002DB6: begin
				q			<=			16'h0741;
		end
		32'h00002DB8: begin
				q			<=			16'h0113;
		end
		32'h00002DBA: begin
				q			<=			16'h0A01;
		end
		32'h00002DBC: begin
				q			<=			16'h8067;
		end
		32'h00002DBE: begin
				q			<=			16'h0000;
		end
		32'h00002DC0: begin
				q			<=			16'h0793;
		end
		32'h00002DC2: begin
				q			<=			16'h2080;
		end
		32'h00002DC4: begin
				q			<=			16'h1A23;
		end
		32'h00002DC6: begin
				q			<=			16'h00F1;
		end
		32'h00002DC8: begin
				q			<=			16'h2423;
		end
		32'h00002DCA: begin
				q			<=			16'h00A1;
		end
		32'h00002DCC: begin
				q			<=			16'h2C23;
		end
		32'h00002DCE: begin
				q			<=			16'h00A1;
		end
		32'h00002DD0: begin
				q			<=			16'h0793;
		end
		32'h00002DD2: begin
				q			<=			16'h0000;
		end
		32'h00002DD4: begin
				q			<=			16'h8463;
		end
		32'h00002DD6: begin
				q			<=			16'h0005;
		end
		32'h00002DD8: begin
				q			<=			16'h8793;
		end
		32'h00002DDA: begin
				q			<=			16'hFFF5;
		end
		32'h00002DDC: begin
				q			<=			16'h2823;
		end
		32'h00002DDE: begin
				q			<=			16'h00F1;
		end
		32'h00002DE0: begin
				q			<=			16'h2E23;
		end
		32'h00002DE2: begin
				q			<=			16'h00F1;
		end
		32'h00002DE4: begin
				q			<=			16'h0693;
		end
		32'h00002DE6: begin
				q			<=			16'h08C1;
		end
		32'h00002DE8: begin
				q			<=			16'h0793;
		end
		32'h00002DEA: begin
				q			<=			16'hFFF0;
		end
		32'h00002DEC: begin
				q			<=			16'h8413;
		end
		32'h00002DEE: begin
				q			<=			16'h0005;
		end
		32'h00002DF0: begin
				q			<=			16'h8513;
		end
		32'h00002DF2: begin
				q			<=			16'h0004;
		end
		32'h00002DF4: begin
				q			<=			16'h0593;
		end
		32'h00002DF6: begin
				q			<=			16'h0081;
		end
		32'h00002DF8: begin
				q			<=			16'h1B23;
		end
		32'h00002DFA: begin
				q			<=			16'h00F1;
		end
		32'h00002DFC: begin
				q			<=			16'h2223;
		end
		32'h00002DFE: begin
				q			<=			16'h00D1;
		end
		32'h00002E00: begin
				q			<=			16'h0097;
		end
		32'h00002E02: begin
				q			<=			16'h0000;
		end
		32'h00002E04: begin
				q			<=			16'h80E7;
		end
		32'h00002E06: begin
				q			<=			16'h0D80;
		end
		32'h00002E08: begin
				q			<=			16'h0793;
		end
		32'h00002E0A: begin
				q			<=			16'hFFF0;
		end
		32'h00002E0C: begin
				q			<=			16'h5663;
		end
		32'h00002E0E: begin
				q			<=			16'h00F5;
		end
		32'h00002E10: begin
				q			<=			16'h0793;
		end
		32'h00002E12: begin
				q			<=			16'h08B0;
		end
		32'h00002E14: begin
				q			<=			16'hA023;
		end
		32'h00002E16: begin
				q			<=			16'h00F4;
		end
		32'h00002E18: begin
				q			<=			16'h0AE3;
		end
		32'h00002E1A: begin
				q			<=			16'hF804;
		end
		32'h00002E1C: begin
				q			<=			16'h2783;
		end
		32'h00002E1E: begin
				q			<=			16'h0081;
		end
		32'h00002E20: begin
				q			<=			16'h8023;
		end
		32'h00002E22: begin
				q			<=			16'h0007;
		end
		32'h00002E24: begin
				q			<=			16'hF06F;
		end
		32'h00002E26: begin
				q			<=			16'hF89F;
		end
		32'h00002E28: begin
				q			<=			16'h0000;
		end
		32'h00002E2A: begin
				q			<=			16'h0000;
		end
		32'h00002E2C: begin
				q			<=			16'h0793;
		end
		32'h00002E2E: begin
				q			<=			16'h0005;
		end
		32'h00002E30: begin
				q			<=			16'h8793;
		end
		32'h00002E32: begin
				q			<=			16'h0017;
		end
		32'h00002E34: begin
				q			<=			16'hC703;
		end
		32'h00002E36: begin
				q			<=			16'hFFF7;
		end
		32'h00002E38: begin
				q			<=			16'h1CE3;
		end
		32'h00002E3A: begin
				q			<=			16'hFE07;
		end
		32'h00002E3C: begin
				q			<=			16'h8533;
		end
		32'h00002E3E: begin
				q			<=			16'h40A7;
		end
		32'h00002E40: begin
				q			<=			16'h0513;
		end
		32'h00002E42: begin
				q			<=			16'hFFF5;
		end
		32'h00002E44: begin
				q			<=			16'h8067;
		end
		32'h00002E46: begin
				q			<=			16'h0000;
		end
		32'h00002E48: begin
				q			<=			16'h0000;
		end
		32'h00002E4A: begin
				q			<=			16'h0000;
		end
		32'h00002E4C: begin
				q			<=			16'h0A63;
		end
		32'h00002E4E: begin
				q			<=			16'h0206;
		end
		32'h00002E50: begin
				q			<=			16'h0713;
		end
		32'h00002E52: begin
				q			<=			16'h0015;
		end
		32'h00002E54: begin
				q			<=			16'h0533;
		end
		32'h00002E56: begin
				q			<=			16'h00C5;
		end
		32'h00002E58: begin
				q			<=			16'h4783;
		end
		32'h00002E5A: begin
				q			<=			16'hFFF7;
		end
		32'h00002E5C: begin
				q			<=			16'hC683;
		end
		32'h00002E5E: begin
				q			<=			16'h0005;
		end
		32'h00002E60: begin
				q			<=			16'h8663;
		end
		32'h00002E62: begin
				q			<=			16'h00D7;
		end
		32'h00002E64: begin
				q			<=			16'h8533;
		end
		32'h00002E66: begin
				q			<=			16'h40D7;
		end
		32'h00002E68: begin
				q			<=			16'h8067;
		end
		32'h00002E6A: begin
				q			<=			16'h0000;
		end
		32'h00002E6C: begin
				q			<=			16'h0CE3;
		end
		32'h00002E6E: begin
				q			<=			16'hFEA7;
		end
		32'h00002E70: begin
				q			<=			16'h0713;
		end
		32'h00002E72: begin
				q			<=			16'h0017;
		end
		32'h00002E74: begin
				q			<=			16'h88E3;
		end
		32'h00002E76: begin
				q			<=			16'hFE07;
		end
		32'h00002E78: begin
				q			<=			16'h8593;
		end
		32'h00002E7A: begin
				q			<=			16'h0015;
		end
		32'h00002E7C: begin
				q			<=			16'hF06F;
		end
		32'h00002E7E: begin
				q			<=			16'hFDDF;
		end
		32'h00002E80: begin
				q			<=			16'h0513;
		end
		32'h00002E82: begin
				q			<=			16'h0000;
		end
		32'h00002E84: begin
				q			<=			16'h8067;
		end
		32'h00002E86: begin
				q			<=			16'h0000;
		end
		32'h00002E88: begin
				q			<=			16'h0000;
		end
		32'h00002E8A: begin
				q			<=			16'h0000;
		end
		32'h00002E8C: begin
				q			<=			16'h0713;
		end
		32'h00002E8E: begin
				q			<=			16'h0005;
		end
		32'h00002E90: begin
				q			<=			16'h1463;
		end
		32'h00002E92: begin
				q			<=			16'h0006;
		end
		32'h00002E94: begin
				q			<=			16'h8067;
		end
		32'h00002E96: begin
				q			<=			16'h0000;
		end
		32'h00002E98: begin
				q			<=			16'h8593;
		end
		32'h00002E9A: begin
				q			<=			16'h0015;
		end
		32'h00002E9C: begin
				q			<=			16'hC683;
		end
		32'h00002E9E: begin
				q			<=			16'hFFF5;
		end
		32'h00002EA0: begin
				q			<=			16'h0793;
		end
		32'h00002EA2: begin
				q			<=			16'h0017;
		end
		32'h00002EA4: begin
				q			<=			16'h0813;
		end
		32'h00002EA6: begin
				q			<=			16'hFFF6;
		end
		32'h00002EA8: begin
				q			<=			16'h8FA3;
		end
		32'h00002EAA: begin
				q			<=			16'hFED7;
		end
		32'h00002EAC: begin
				q			<=			16'h9863;
		end
		32'h00002EAE: begin
				q			<=			16'h0006;
		end
		32'h00002EB0: begin
				q			<=			16'h0733;
		end
		32'h00002EB2: begin
				q			<=			16'h00C7;
		end
		32'h00002EB4: begin
				q			<=			16'h9A63;
		end
		32'h00002EB6: begin
				q			<=			16'h00E7;
		end
		32'h00002EB8: begin
				q			<=			16'h8067;
		end
		32'h00002EBA: begin
				q			<=			16'h0000;
		end
		32'h00002EBC: begin
				q			<=			16'h8713;
		end
		32'h00002EBE: begin
				q			<=			16'h0007;
		end
		32'h00002EC0: begin
				q			<=			16'h0613;
		end
		32'h00002EC2: begin
				q			<=			16'h0008;
		end
		32'h00002EC4: begin
				q			<=			16'hF06F;
		end
		32'h00002EC6: begin
				q			<=			16'hFCDF;
		end
		32'h00002EC8: begin
				q			<=			16'h8793;
		end
		32'h00002ECA: begin
				q			<=			16'h0017;
		end
		32'h00002ECC: begin
				q			<=			16'h8FA3;
		end
		32'h00002ECE: begin
				q			<=			16'hFE07;
		end
		32'h00002ED0: begin
				q			<=			16'hF06F;
		end
		32'h00002ED2: begin
				q			<=			16'hFE5F;
		end
		32'h00002ED4: begin
				q			<=			16'h0000;
		end
		32'h00002ED6: begin
				q			<=			16'h0000;
		end
		32'h00002ED8: begin
				q			<=			16'h0113;
		end
		32'h00002EDA: begin
				q			<=			16'hE301;
		end
		32'h00002EDC: begin
				q			<=			16'h2623;
		end
		32'h00002EDE: begin
				q			<=			16'h1C11;
		end
		32'h00002EE0: begin
				q			<=			16'h2223;
		end
		32'h00002EE2: begin
				q			<=			16'h1C91;
		end
		32'h00002EE4: begin
				q			<=			16'h2023;
		end
		32'h00002EE6: begin
				q			<=			16'h1D21;
		end
		32'h00002EE8: begin
				q			<=			16'h2E23;
		end
		32'h00002EEA: begin
				q			<=			16'h1B31;
		end
		32'h00002EEC: begin
				q			<=			16'h2A23;
		end
		32'h00002EEE: begin
				q			<=			16'h1B51;
		end
		32'h00002EF0: begin
				q			<=			16'h8993;
		end
		32'h00002EF2: begin
				q			<=			16'h0005;
		end
		32'h00002EF4: begin
				q			<=			16'h0493;
		end
		32'h00002EF6: begin
				q			<=			16'h0006;
		end
		32'h00002EF8: begin
				q			<=			16'h8A93;
		end
		32'h00002EFA: begin
				q			<=			16'h0006;
		end
		32'h00002EFC: begin
				q			<=			16'h2423;
		end
		32'h00002EFE: begin
				q			<=			16'h1C81;
		end
		32'h00002F00: begin
				q			<=			16'h2C23;
		end
		32'h00002F02: begin
				q			<=			16'h1B41;
		end
		32'h00002F04: begin
				q			<=			16'h2823;
		end
		32'h00002F06: begin
				q			<=			16'h1B61;
		end
		32'h00002F08: begin
				q			<=			16'h2623;
		end
		32'h00002F0A: begin
				q			<=			16'h1B71;
		end
		32'h00002F0C: begin
				q			<=			16'h2423;
		end
		32'h00002F0E: begin
				q			<=			16'h1B81;
		end
		32'h00002F10: begin
				q			<=			16'h2223;
		end
		32'h00002F12: begin
				q			<=			16'h1B91;
		end
		32'h00002F14: begin
				q			<=			16'h2023;
		end
		32'h00002F16: begin
				q			<=			16'h1BA1;
		end
		32'h00002F18: begin
				q			<=			16'h2E23;
		end
		32'h00002F1A: begin
				q			<=			16'h19B1;
		end
		32'h00002F1C: begin
				q			<=			16'h0913;
		end
		32'h00002F1E: begin
				q			<=			16'h0005;
		end
		32'h00002F20: begin
				q			<=			16'h4097;
		end
		32'h00002F22: begin
				q			<=			16'h0000;
		end
		32'h00002F24: begin
				q			<=			16'h80E7;
		end
		32'h00002F26: begin
				q			<=			16'h4340;
		end
		32'h00002F28: begin
				q			<=			16'h2783;
		end
		32'h00002F2A: begin
				q			<=			16'h0005;
		end
		32'h00002F2C: begin
				q			<=			16'h8513;
		end
		32'h00002F2E: begin
				q			<=			16'h0007;
		end
		32'h00002F30: begin
				q			<=			16'h2423;
		end
		32'h00002F32: begin
				q			<=			16'h02F1;
		end
		32'h00002F34: begin
				q			<=			16'hF0EF;
		end
		32'h00002F36: begin
				q			<=			16'hEF9F;
		end
		32'h00002F38: begin
				q			<=			16'hD783;
		end
		32'h00002F3A: begin
				q			<=			16'h00C9;
		end
		32'h00002F3C: begin
				q			<=			16'h2A23;
		end
		32'h00002F3E: begin
				q			<=			16'h00A1;
		end
		32'h00002F40: begin
				q			<=			16'h2823;
		end
		32'h00002F42: begin
				q			<=			16'h0C01;
		end
		32'h00002F44: begin
				q			<=			16'h2A23;
		end
		32'h00002F46: begin
				q			<=			16'h0C01;
		end
		32'h00002F48: begin
				q			<=			16'h2C23;
		end
		32'h00002F4A: begin
				q			<=			16'h0C01;
		end
		32'h00002F4C: begin
				q			<=			16'h2E23;
		end
		32'h00002F4E: begin
				q			<=			16'h0C01;
		end
		32'h00002F50: begin
				q			<=			16'hF793;
		end
		32'h00002F52: begin
				q			<=			16'h0807;
		end
		32'h00002F54: begin
				q			<=			16'h8063;
		end
		32'h00002F56: begin
				q			<=			16'h0407;
		end
		32'h00002F58: begin
				q			<=			16'hA783;
		end
		32'h00002F5A: begin
				q			<=			16'h0109;
		end
		32'h00002F5C: begin
				q			<=			16'h9C63;
		end
		32'h00002F5E: begin
				q			<=			16'h0207;
		end
		32'h00002F60: begin
				q			<=			16'h0593;
		end
		32'h00002F62: begin
				q			<=			16'h0400;
		end
		32'h00002F64: begin
				q			<=			16'h0513;
		end
		32'h00002F66: begin
				q			<=			16'h0009;
		end
		32'h00002F68: begin
				q			<=			16'h40EF;
		end
		32'h00002F6A: begin
				q			<=			16'h4380;
		end
		32'h00002F6C: begin
				q			<=			16'hA023;
		end
		32'h00002F6E: begin
				q			<=			16'h00A9;
		end
		32'h00002F70: begin
				q			<=			16'hA823;
		end
		32'h00002F72: begin
				q			<=			16'h00A9;
		end
		32'h00002F74: begin
				q			<=			16'h1C63;
		end
		32'h00002F76: begin
				q			<=			16'h0005;
		end
		32'h00002F78: begin
				q			<=			16'h0793;
		end
		32'h00002F7A: begin
				q			<=			16'h00C0;
		end
		32'h00002F7C: begin
				q			<=			16'h2023;
		end
		32'h00002F7E: begin
				q			<=			16'h00F9;
		end
		32'h00002F80: begin
				q			<=			16'h0793;
		end
		32'h00002F82: begin
				q			<=			16'hFFF0;
		end
		32'h00002F84: begin
				q			<=			16'h2C23;
		end
		32'h00002F86: begin
				q			<=			16'h00F1;
		end
		32'h00002F88: begin
				q			<=			16'h006F;
		end
		32'h00002F8A: begin
				q			<=			16'h5840;
		end
		32'h00002F8C: begin
				q			<=			16'h0793;
		end
		32'h00002F8E: begin
				q			<=			16'h0400;
		end
		32'h00002F90: begin
				q			<=			16'hAA23;
		end
		32'h00002F92: begin
				q			<=			16'h00F9;
		end
		32'h00002F94: begin
				q			<=			16'h0893;
		end
		32'h00002F96: begin
				q			<=			16'h0EC1;
		end
		32'h00002F98: begin
				q			<=			16'h2223;
		end
		32'h00002F9A: begin
				q			<=			16'h0D11;
		end
		32'h00002F9C: begin
				q			<=			16'h2623;
		end
		32'h00002F9E: begin
				q			<=			16'h0C01;
		end
		32'h00002FA0: begin
				q			<=			16'h2423;
		end
		32'h00002FA2: begin
				q			<=			16'h0C01;
		end
		32'h00002FA4: begin
				q			<=			16'h0A13;
		end
		32'h00002FA6: begin
				q			<=			16'h0000;
		end
		32'h00002FA8: begin
				q			<=			16'h2A23;
		end
		32'h00002FAA: begin
				q			<=			16'h0201;
		end
		32'h00002FAC: begin
				q			<=			16'h2823;
		end
		32'h00002FAE: begin
				q			<=			16'h0201;
		end
		32'h00002FB0: begin
				q			<=			16'h2423;
		end
		32'h00002FB2: begin
				q			<=			16'h0001;
		end
		32'h00002FB4: begin
				q			<=			16'h2223;
		end
		32'h00002FB6: begin
				q			<=			16'h0201;
		end
		32'h00002FB8: begin
				q			<=			16'h2623;
		end
		32'h00002FBA: begin
				q			<=			16'h0201;
		end
		32'h00002FBC: begin
				q			<=			16'h2C23;
		end
		32'h00002FBE: begin
				q			<=			16'h0001;
		end
		32'h00002FC0: begin
				q			<=			16'h8413;
		end
		32'h00002FC2: begin
				q			<=			16'h0004;
		end
		32'h00002FC4: begin
				q			<=			16'h0713;
		end
		32'h00002FC6: begin
				q			<=			16'h0250;
		end
		32'h00002FC8: begin
				q			<=			16'h4783;
		end
		32'h00002FCA: begin
				q			<=			16'h0004;
		end
		32'h00002FCC: begin
				q			<=			16'h8463;
		end
		32'h00002FCE: begin
				q			<=			16'h0007;
		end
		32'h00002FD0: begin
				q			<=			16'h9263;
		end
		32'h00002FD2: begin
				q			<=			16'h0CE7;
		end
		32'h00002FD4: begin
				q			<=			16'h0B33;
		end
		32'h00002FD6: begin
				q			<=			16'h4094;
		end
		32'h00002FD8: begin
				q			<=			16'h0A63;
		end
		32'h00002FDA: begin
				q			<=			16'h040B;
		end
		32'h00002FDC: begin
				q			<=			16'h2783;
		end
		32'h00002FDE: begin
				q			<=			16'h0CC1;
		end
		32'h00002FE0: begin
				q			<=			16'hA023;
		end
		32'h00002FE2: begin
				q			<=			16'h0098;
		end
		32'h00002FE4: begin
				q			<=			16'hA223;
		end
		32'h00002FE6: begin
				q			<=			16'h0168;
		end
		32'h00002FE8: begin
				q			<=			16'h87B3;
		end
		32'h00002FEA: begin
				q			<=			16'h0167;
		end
		32'h00002FEC: begin
				q			<=			16'h2623;
		end
		32'h00002FEE: begin
				q			<=			16'h0CF1;
		end
		32'h00002FF0: begin
				q			<=			16'h2783;
		end
		32'h00002FF2: begin
				q			<=			16'h0C81;
		end
		32'h00002FF4: begin
				q			<=			16'h0713;
		end
		32'h00002FF6: begin
				q			<=			16'h0070;
		end
		32'h00002FF8: begin
				q			<=			16'h8893;
		end
		32'h00002FFA: begin
				q			<=			16'h0088;
		end
		32'h00002FFC: begin
				q			<=			16'h8793;
		end
		32'h00002FFE: begin
				q			<=			16'h0017;
		end
		32'h00003000: begin
				q			<=			16'h2423;
		end
		32'h00003002: begin
				q			<=			16'h0CF1;
		end
		32'h00003004: begin
				q			<=			16'h5E63;
		end
		32'h00003006: begin
				q			<=			16'h00F7;
		end
		32'h00003008: begin
				q			<=			16'h0613;
		end
		32'h0000300A: begin
				q			<=			16'h0C41;
		end
		32'h0000300C: begin
				q			<=			16'h8593;
		end
		32'h0000300E: begin
				q			<=			16'h0009;
		end
		32'h00003010: begin
				q			<=			16'h0513;
		end
		32'h00003012: begin
				q			<=			16'h0009;
		end
		32'h00003014: begin
				q			<=			16'h50EF;
		end
		32'h00003016: begin
				q			<=			16'h3490;
		end
		32'h00003018: begin
				q			<=			16'h1463;
		end
		32'h0000301A: begin
				q			<=			16'h4E05;
		end
		32'h0000301C: begin
				q			<=			16'h0893;
		end
		32'h0000301E: begin
				q			<=			16'h0EC1;
		end
		32'h00003020: begin
				q			<=			16'h2783;
		end
		32'h00003022: begin
				q			<=			16'h0181;
		end
		32'h00003024: begin
				q			<=			16'h87B3;
		end
		32'h00003026: begin
				q			<=			16'h0167;
		end
		32'h00003028: begin
				q			<=			16'h2C23;
		end
		32'h0000302A: begin
				q			<=			16'h00F1;
		end
		32'h0000302C: begin
				q			<=			16'h4783;
		end
		32'h0000302E: begin
				q			<=			16'h0004;
		end
		32'h00003030: begin
				q			<=			16'h9463;
		end
		32'h00003032: begin
				q			<=			16'h0007;
		end
		32'h00003034: begin
				q			<=			16'h106F;
		end
		32'h00003036: begin
				q			<=			16'h5E90;
		end
		32'h00003038: begin
				q			<=			16'h0793;
		end
		32'h0000303A: begin
				q			<=			16'h0014;
		end
		32'h0000303C: begin
				q			<=			16'h2823;
		end
		32'h0000303E: begin
				q			<=			16'h00F1;
		end
		32'h00003040: begin
				q			<=			16'h03A3;
		end
		32'h00003042: begin
				q			<=			16'h0A01;
		end
		32'h00003044: begin
				q			<=			16'h0B13;
		end
		32'h00003046: begin
				q			<=			16'hFFF0;
		end
		32'h00003048: begin
				q			<=			16'h2E23;
		end
		32'h0000304A: begin
				q			<=			16'h0001;
		end
		32'h0000304C: begin
				q			<=			16'h0413;
		end
		32'h0000304E: begin
				q			<=			16'h0000;
		end
		32'h00003050: begin
				q			<=			16'h0B93;
		end
		32'h00003052: begin
				q			<=			16'h0090;
		end
		32'h00003054: begin
				q			<=			16'h0693;
		end
		32'h00003056: begin
				q			<=			16'h05A0;
		end
		32'h00003058: begin
				q			<=			16'h0613;
		end
		32'h0000305A: begin
				q			<=			16'h02A0;
		end
		32'h0000305C: begin
				q			<=			16'h2783;
		end
		32'h0000305E: begin
				q			<=			16'h0101;
		end
		32'h00003060: begin
				q			<=			16'hCD03;
		end
		32'h00003062: begin
				q			<=			16'h0007;
		end
		32'h00003064: begin
				q			<=			16'h8793;
		end
		32'h00003066: begin
				q			<=			16'h0017;
		end
		32'h00003068: begin
				q			<=			16'h2823;
		end
		32'h0000306A: begin
				q			<=			16'h00F1;
		end
		32'h0000306C: begin
				q			<=			16'h0793;
		end
		32'h0000306E: begin
				q			<=			16'hFE0D;
		end
		32'h00003070: begin
				q			<=			16'hF463;
		end
		32'h00003072: begin
				q			<=			16'h00F6;
		end
		32'h00003074: begin
				q			<=			16'h106F;
		end
		32'h00003076: begin
				q			<=			16'h2A40;
		end
		32'h00003078: begin
				q			<=			16'hC717;
		end
		32'h0000307A: begin
				q			<=			16'h0000;
		end
		32'h0000307C: begin
				q			<=			16'h0713;
		end
		32'h0000307E: begin
				q			<=			16'h0A87;
		end
		32'h00003080: begin
				q			<=			16'h9793;
		end
		32'h00003082: begin
				q			<=			16'h0027;
		end
		32'h00003084: begin
				q			<=			16'h87B3;
		end
		32'h00003086: begin
				q			<=			16'h00E7;
		end
		32'h00003088: begin
				q			<=			16'hA783;
		end
		32'h0000308A: begin
				q			<=			16'h0007;
		end
		32'h0000308C: begin
				q			<=			16'h87B3;
		end
		32'h0000308E: begin
				q			<=			16'h00E7;
		end
		32'h00003090: begin
				q			<=			16'h8067;
		end
		32'h00003092: begin
				q			<=			16'h0007;
		end
		32'h00003094: begin
				q			<=			16'h0413;
		end
		32'h00003096: begin
				q			<=			16'h0014;
		end
		32'h00003098: begin
				q			<=			16'hF06F;
		end
		32'h0000309A: begin
				q			<=			16'hF31F;
		end
		32'h0000309C: begin
				q			<=			16'hD797;
		end
		32'h0000309E: begin
				q			<=			16'h0000;
		end
		32'h000030A0: begin
				q			<=			16'h8793;
		end
		32'h000030A2: begin
				q			<=			16'hCFC7;
		end
		32'h000030A4: begin
				q			<=			16'h2A23;
		end
		32'h000030A6: begin
				q			<=			16'h02F1;
		end
		32'h000030A8: begin
				q			<=			16'h7793;
		end
		32'h000030AA: begin
				q			<=			16'h0204;
		end
		32'h000030AC: begin
				q			<=			16'h9463;
		end
		32'h000030AE: begin
				q			<=			16'h0007;
		end
		32'h000030B0: begin
				q			<=			16'h106F;
		end
		32'h000030B2: begin
				q			<=			16'h0840;
		end
		32'h000030B4: begin
				q			<=			16'h8A93;
		end
		32'h000030B6: begin
				q			<=			16'h007A;
		end
		32'h000030B8: begin
				q			<=			16'hFA93;
		end
		32'h000030BA: begin
				q			<=			16'hFF8A;
		end
		32'h000030BC: begin
				q			<=			16'hAC03;
		end
		32'h000030BE: begin
				q			<=			16'h000A;
		end
		32'h000030C0: begin
				q			<=			16'hAC83;
		end
		32'h000030C2: begin
				q			<=			16'h004A;
		end
		32'h000030C4: begin
				q			<=			16'h8793;
		end
		32'h000030C6: begin
				q			<=			16'h008A;
		end
		32'h000030C8: begin
				q			<=			16'h2623;
		end
		32'h000030CA: begin
				q			<=			16'h00F1;
		end
		32'h000030CC: begin
				q			<=			16'h7793;
		end
		32'h000030CE: begin
				q			<=			16'h0014;
		end
		32'h000030D0: begin
				q			<=			16'h8E63;
		end
		32'h000030D2: begin
				q			<=			16'h0007;
		end
		32'h000030D4: begin
				q			<=			16'h67B3;
		end
		32'h000030D6: begin
				q			<=			16'h019C;
		end
		32'h000030D8: begin
				q			<=			16'h8A63;
		end
		32'h000030DA: begin
				q			<=			16'h0007;
		end
		32'h000030DC: begin
				q			<=			16'h0793;
		end
		32'h000030DE: begin
				q			<=			16'h0300;
		end
		32'h000030E0: begin
				q			<=			16'h0423;
		end
		32'h000030E2: begin
				q			<=			16'h0AF1;
		end
		32'h000030E4: begin
				q			<=			16'h04A3;
		end
		32'h000030E6: begin
				q			<=			16'h0BA1;
		end
		32'h000030E8: begin
				q			<=			16'h6413;
		end
		32'h000030EA: begin
				q			<=			16'h0024;
		end
		32'h000030EC: begin
				q			<=			16'h7413;
		end
		32'h000030EE: begin
				q			<=			16'hBFF4;
		end
		32'h000030F0: begin
				q			<=			16'h0793;
		end
		32'h000030F2: begin
				q			<=			16'h0020;
		end
		32'h000030F4: begin
				q			<=			16'h006F;
		end
		32'h000030F6: begin
				q			<=			16'h4490;
		end
		32'h000030F8: begin
				q			<=			16'h0513;
		end
		32'h000030FA: begin
				q			<=			16'h0009;
		end
		32'h000030FC: begin
				q			<=			16'h2223;
		end
		32'h000030FE: begin
				q			<=			16'h0111;
		end
		32'h00003100: begin
				q			<=			16'h4097;
		end
		32'h00003102: begin
				q			<=			16'h0000;
		end
		32'h00003104: begin
				q			<=			16'h80E7;
		end
		32'h00003106: begin
				q			<=			16'h2540;
		end
		32'h00003108: begin
				q			<=			16'h2783;
		end
		32'h0000310A: begin
				q			<=			16'h0045;
		end
		32'h0000310C: begin
				q			<=			16'h8513;
		end
		32'h0000310E: begin
				q			<=			16'h0007;
		end
		32'h00003110: begin
				q			<=			16'h2623;
		end
		32'h00003112: begin
				q			<=			16'h02F1;
		end
		32'h00003114: begin
				q			<=			16'hF0EF;
		end
		32'h00003116: begin
				q			<=			16'hD19F;
		end
		32'h00003118: begin
				q			<=			16'h2223;
		end
		32'h0000311A: begin
				q			<=			16'h02A1;
		end
		32'h0000311C: begin
				q			<=			16'h0513;
		end
		32'h0000311E: begin
				q			<=			16'h0009;
		end
		32'h00003120: begin
				q			<=			16'h4097;
		end
		32'h00003122: begin
				q			<=			16'h0000;
		end
		32'h00003124: begin
				q			<=			16'h80E7;
		end
		32'h00003126: begin
				q			<=			16'h2340;
		end
		32'h00003128: begin
				q			<=			16'h2783;
		end
		32'h0000312A: begin
				q			<=			16'h0085;
		end
		32'h0000312C: begin
				q			<=			16'h2883;
		end
		32'h0000312E: begin
				q			<=			16'h0041;
		end
		32'h00003130: begin
				q			<=			16'h2423;
		end
		32'h00003132: begin
				q			<=			16'h00F1;
		end
		32'h00003134: begin
				q			<=			16'h2783;
		end
		32'h00003136: begin
				q			<=			16'h0241;
		end
		32'h00003138: begin
				q			<=			16'h8EE3;
		end
		32'h0000313A: begin
				q			<=			16'hF007;
		end
		32'h0000313C: begin
				q			<=			16'h2783;
		end
		32'h0000313E: begin
				q			<=			16'h0081;
		end
		32'h00003140: begin
				q			<=			16'h8AE3;
		end
		32'h00003142: begin
				q			<=			16'hF007;
		end
		32'h00003144: begin
				q			<=			16'hC783;
		end
		32'h00003146: begin
				q			<=			16'h0007;
		end
		32'h00003148: begin
				q			<=			16'h86E3;
		end
		32'h0000314A: begin
				q			<=			16'hF007;
		end
		32'h0000314C: begin
				q			<=			16'h6413;
		end
		32'h0000314E: begin
				q			<=			16'h4004;
		end
		32'h00003150: begin
				q			<=			16'hF06F;
		end
		32'h00003152: begin
				q			<=			16'hF05F;
		end
		32'h00003154: begin
				q			<=			16'h4783;
		end
		32'h00003156: begin
				q			<=			16'h0A71;
		end
		32'h00003158: begin
				q			<=			16'h9EE3;
		end
		32'h0000315A: begin
				q			<=			16'hEE07;
		end
		32'h0000315C: begin
				q			<=			16'h0793;
		end
		32'h0000315E: begin
				q			<=			16'h0200;
		end
		32'h00003160: begin
				q			<=			16'h03A3;
		end
		32'h00003162: begin
				q			<=			16'h0AF1;
		end
		32'h00003164: begin
				q			<=			16'hF06F;
		end
		32'h00003166: begin
				q			<=			16'hEF1F;
		end
		32'h00003168: begin
				q			<=			16'h6413;
		end
		32'h0000316A: begin
				q			<=			16'h0014;
		end
		32'h0000316C: begin
				q			<=			16'hF06F;
		end
		32'h0000316E: begin
				q			<=			16'hEE9F;
		end
		32'h00003170: begin
				q			<=			16'hA783;
		end
		32'h00003172: begin
				q			<=			16'h000A;
		end
		32'h00003174: begin
				q			<=			16'h8A93;
		end
		32'h00003176: begin
				q			<=			16'h004A;
		end
		32'h00003178: begin
				q			<=			16'h2E23;
		end
		32'h0000317A: begin
				q			<=			16'h00F1;
		end
		32'h0000317C: begin
				q			<=			16'hDCE3;
		end
		32'h0000317E: begin
				q			<=			16'hEC07;
		end
		32'h00003180: begin
				q			<=			16'h07B3;
		end
		32'h00003182: begin
				q			<=			16'h40F0;
		end
		32'h00003184: begin
				q			<=			16'h2E23;
		end
		32'h00003186: begin
				q			<=			16'h00F1;
		end
		32'h00003188: begin
				q			<=			16'h6413;
		end
		32'h0000318A: begin
				q			<=			16'h0044;
		end
		32'h0000318C: begin
				q			<=			16'hF06F;
		end
		32'h0000318E: begin
				q			<=			16'hEC9F;
		end
		32'h00003190: begin
				q			<=			16'h0793;
		end
		32'h00003192: begin
				q			<=			16'h02B0;
		end
		32'h00003194: begin
				q			<=			16'hF06F;
		end
		32'h00003196: begin
				q			<=			16'hFCDF;
		end
		32'h00003198: begin
				q			<=			16'h2703;
		end
		32'h0000319A: begin
				q			<=			16'h0101;
		end
		32'h0000319C: begin
				q			<=			16'h2783;
		end
		32'h0000319E: begin
				q			<=			16'h0101;
		end
		32'h000031A0: begin
				q			<=			16'h4D03;
		end
		32'h000031A2: begin
				q			<=			16'h0007;
		end
		32'h000031A4: begin
				q			<=			16'h8793;
		end
		32'h000031A6: begin
				q			<=			16'h0017;
		end
		32'h000031A8: begin
				q			<=			16'h1063;
		end
		32'h000031AA: begin
				q			<=			16'h04CD;
		end
		32'h000031AC: begin
				q			<=			16'hAB03;
		end
		32'h000031AE: begin
				q			<=			16'h000A;
		end
		32'h000031B0: begin
				q			<=			16'h8713;
		end
		32'h000031B2: begin
				q			<=			16'h004A;
		end
		32'h000031B4: begin
				q			<=			16'h5463;
		end
		32'h000031B6: begin
				q			<=			16'h000B;
		end
		32'h000031B8: begin
				q			<=			16'h0B13;
		end
		32'h000031BA: begin
				q			<=			16'hFFF0;
		end
		32'h000031BC: begin
				q			<=			16'h0A93;
		end
		32'h000031BE: begin
				q			<=			16'h0007;
		end
		32'h000031C0: begin
				q			<=			16'h2823;
		end
		32'h000031C2: begin
				q			<=			16'h00F1;
		end
		32'h000031C4: begin
				q			<=			16'hF06F;
		end
		32'h000031C6: begin
				q			<=			16'hE91F;
		end
		32'h000031C8: begin
				q			<=			16'h0593;
		end
		32'h000031CA: begin
				q			<=			16'h00A0;
		end
		32'h000031CC: begin
				q			<=			16'h0333;
		end
		32'h000031CE: begin
				q			<=			16'h02BB;
		end
		32'h000031D0: begin
				q			<=			16'h8793;
		end
		32'h000031D2: begin
				q			<=			16'h0017;
		end
		32'h000031D4: begin
				q			<=			16'hCD03;
		end
		32'h000031D6: begin
				q			<=			16'hFFF7;
		end
		32'h000031D8: begin
				q			<=			16'h0B33;
		end
		32'h000031DA: begin
				q			<=			16'h00E3;
		end
		32'h000031DC: begin
				q			<=			16'h0713;
		end
		32'h000031DE: begin
				q			<=			16'hFD0D;
		end
		32'h000031E0: begin
				q			<=			16'hF4E3;
		end
		32'h000031E2: begin
				q			<=			16'hFEEB;
		end
		32'h000031E4: begin
				q			<=			16'hF06F;
		end
		32'h000031E6: begin
				q			<=			16'hE85F;
		end
		32'h000031E8: begin
				q			<=			16'h0B13;
		end
		32'h000031EA: begin
				q			<=			16'h0000;
		end
		32'h000031EC: begin
				q			<=			16'hF06F;
		end
		32'h000031EE: begin
				q			<=			16'hFF1F;
		end
		32'h000031F0: begin
				q			<=			16'h6413;
		end
		32'h000031F2: begin
				q			<=			16'h0804;
		end
		32'h000031F4: begin
				q			<=			16'hF06F;
		end
		32'h000031F6: begin
				q			<=			16'hE61F;
		end
		32'h000031F8: begin
				q			<=			16'h2783;
		end
		32'h000031FA: begin
				q			<=			16'h0101;
		end
		32'h000031FC: begin
				q			<=			16'h2E23;
		end
		32'h000031FE: begin
				q			<=			16'h0001;
		end
		32'h00003200: begin
				q			<=			16'h2703;
		end
		32'h00003202: begin
				q			<=			16'h01C1;
		end
		32'h00003204: begin
				q			<=			16'h0593;
		end
		32'h00003206: begin
				q			<=			16'h00A0;
		end
		32'h00003208: begin
				q			<=			16'h0D13;
		end
		32'h0000320A: begin
				q			<=			16'hFD0D;
		end
		32'h0000320C: begin
				q			<=			16'h0733;
		end
		32'h0000320E: begin
				q			<=			16'h02B7;
		end
		32'h00003210: begin
				q			<=			16'h8793;
		end
		32'h00003212: begin
				q			<=			16'h0017;
		end
		32'h00003214: begin
				q			<=			16'h0733;
		end
		32'h00003216: begin
				q			<=			16'h00ED;
		end
		32'h00003218: begin
				q			<=			16'hCD03;
		end
		32'h0000321A: begin
				q			<=			16'hFFF7;
		end
		32'h0000321C: begin
				q			<=			16'h2E23;
		end
		32'h0000321E: begin
				q			<=			16'h00E1;
		end
		32'h00003220: begin
				q			<=			16'h0713;
		end
		32'h00003222: begin
				q			<=			16'hFD0D;
		end
		32'h00003224: begin
				q			<=			16'hFEE3;
		end
		32'h00003226: begin
				q			<=			16'hFCEB;
		end
		32'h00003228: begin
				q			<=			16'hF06F;
		end
		32'h0000322A: begin
				q			<=			16'hE41F;
		end
		32'h0000322C: begin
				q			<=			16'h6413;
		end
		32'h0000322E: begin
				q			<=			16'h0084;
		end
		32'h00003230: begin
				q			<=			16'hF06F;
		end
		32'h00003232: begin
				q			<=			16'hE25F;
		end
		32'h00003234: begin
				q			<=			16'h2783;
		end
		32'h00003236: begin
				q			<=			16'h0101;
		end
		32'h00003238: begin
				q			<=			16'hC703;
		end
		32'h0000323A: begin
				q			<=			16'h0007;
		end
		32'h0000323C: begin
				q			<=			16'h0793;
		end
		32'h0000323E: begin
				q			<=			16'h0680;
		end
		32'h00003240: begin
				q			<=			16'h1C63;
		end
		32'h00003242: begin
				q			<=			16'h00F7;
		end
		32'h00003244: begin
				q			<=			16'h2783;
		end
		32'h00003246: begin
				q			<=			16'h0101;
		end
		32'h00003248: begin
				q			<=			16'h6413;
		end
		32'h0000324A: begin
				q			<=			16'h2004;
		end
		32'h0000324C: begin
				q			<=			16'h8793;
		end
		32'h0000324E: begin
				q			<=			16'h0017;
		end
		32'h00003250: begin
				q			<=			16'h2823;
		end
		32'h00003252: begin
				q			<=			16'h00F1;
		end
		32'h00003254: begin
				q			<=			16'hF06F;
		end
		32'h00003256: begin
				q			<=			16'hE01F;
		end
		32'h00003258: begin
				q			<=			16'h6413;
		end
		32'h0000325A: begin
				q			<=			16'h0404;
		end
		32'h0000325C: begin
				q			<=			16'hF06F;
		end
		32'h0000325E: begin
				q			<=			16'hDF9F;
		end
		32'h00003260: begin
				q			<=			16'h2783;
		end
		32'h00003262: begin
				q			<=			16'h0101;
		end
		32'h00003264: begin
				q			<=			16'hC703;
		end
		32'h00003266: begin
				q			<=			16'h0007;
		end
		32'h00003268: begin
				q			<=			16'h0793;
		end
		32'h0000326A: begin
				q			<=			16'h06C0;
		end
		32'h0000326C: begin
				q			<=			16'h1C63;
		end
		32'h0000326E: begin
				q			<=			16'h00F7;
		end
		32'h00003270: begin
				q			<=			16'h2783;
		end
		32'h00003272: begin
				q			<=			16'h0101;
		end
		32'h00003274: begin
				q			<=			16'h8793;
		end
		32'h00003276: begin
				q			<=			16'h0017;
		end
		32'h00003278: begin
				q			<=			16'h2823;
		end
		32'h0000327A: begin
				q			<=			16'h00F1;
		end
		32'h0000327C: begin
				q			<=			16'h6413;
		end
		32'h0000327E: begin
				q			<=			16'h0204;
		end
		32'h00003280: begin
				q			<=			16'hF06F;
		end
		32'h00003282: begin
				q			<=			16'hDD5F;
		end
		32'h00003284: begin
				q			<=			16'h6413;
		end
		32'h00003286: begin
				q			<=			16'h0104;
		end
		32'h00003288: begin
				q			<=			16'hF06F;
		end
		32'h0000328A: begin
				q			<=			16'hDCDF;
		end
		32'h0000328C: begin
				q			<=			16'h8793;
		end
		32'h0000328E: begin
				q			<=			16'h004A;
		end
		32'h00003290: begin
				q			<=			16'h2623;
		end
		32'h00003292: begin
				q			<=			16'h00F1;
		end
		32'h00003294: begin
				q			<=			16'hA783;
		end
		32'h00003296: begin
				q			<=			16'h000A;
		end
		32'h00003298: begin
				q			<=			16'h03A3;
		end
		32'h0000329A: begin
				q			<=			16'h0A01;
		end
		32'h0000329C: begin
				q			<=			16'h0623;
		end
		32'h0000329E: begin
				q			<=			16'h12F1;
		end
		32'h000032A0: begin
				q			<=			16'h2223;
		end
		32'h000032A2: begin
				q			<=			16'h0001;
		end
		32'h000032A4: begin
				q			<=			16'h0B13;
		end
		32'h000032A6: begin
				q			<=			16'h0010;
		end
		32'h000032A8: begin
				q			<=			16'h0D93;
		end
		32'h000032AA: begin
				q			<=			16'h0000;
		end
		32'h000032AC: begin
				q			<=			16'h0C13;
		end
		32'h000032AE: begin
				q			<=			16'h0000;
		end
		32'h000032B0: begin
				q			<=			16'h0B93;
		end
		32'h000032B2: begin
				q			<=			16'h0000;
		end
		32'h000032B4: begin
				q			<=			16'h0C93;
		end
		32'h000032B6: begin
				q			<=			16'h0000;
		end
		32'h000032B8: begin
				q			<=			16'h0493;
		end
		32'h000032BA: begin
				q			<=			16'h12C1;
		end
		32'h000032BC: begin
				q			<=			16'h006F;
		end
		32'h000032BE: begin
				q			<=			16'h3890;
		end
		32'h000032C0: begin
				q			<=			16'h6413;
		end
		32'h000032C2: begin
				q			<=			16'h0104;
		end
		32'h000032C4: begin
				q			<=			16'h7793;
		end
		32'h000032C6: begin
				q			<=			16'h0204;
		end
		32'h000032C8: begin
				q			<=			16'h8E63;
		end
		32'h000032CA: begin
				q			<=			16'h0407;
		end
		32'h000032CC: begin
				q			<=			16'h8A93;
		end
		32'h000032CE: begin
				q			<=			16'h007A;
		end
		32'h000032D0: begin
				q			<=			16'hFA93;
		end
		32'h000032D2: begin
				q			<=			16'hFF8A;
		end
		32'h000032D4: begin
				q			<=			16'hAC03;
		end
		32'h000032D6: begin
				q			<=			16'h000A;
		end
		32'h000032D8: begin
				q			<=			16'hAC83;
		end
		32'h000032DA: begin
				q			<=			16'h004A;
		end
		32'h000032DC: begin
				q			<=			16'h8793;
		end
		32'h000032DE: begin
				q			<=			16'h008A;
		end
		32'h000032E0: begin
				q			<=			16'h2623;
		end
		32'h000032E2: begin
				q			<=			16'h00F1;
		end
		32'h000032E4: begin
				q			<=			16'hDE63;
		end
		32'h000032E6: begin
				q			<=			16'h000C;
		end
		32'h000032E8: begin
				q			<=			16'h0C33;
		end
		32'h000032EA: begin
				q			<=			16'h4180;
		end
		32'h000032EC: begin
				q			<=			16'h37B3;
		end
		32'h000032EE: begin
				q			<=			16'h0180;
		end
		32'h000032F0: begin
				q			<=			16'h0CB3;
		end
		32'h000032F2: begin
				q			<=			16'h4190;
		end
		32'h000032F4: begin
				q			<=			16'h8CB3;
		end
		32'h000032F6: begin
				q			<=			16'h40FC;
		end
		32'h000032F8: begin
				q			<=			16'h0793;
		end
		32'h000032FA: begin
				q			<=			16'h02D0;
		end
		32'h000032FC: begin
				q			<=			16'h03A3;
		end
		32'h000032FE: begin
				q			<=			16'h0AF1;
		end
		32'h00003300: begin
				q			<=			16'h0793;
		end
		32'h00003302: begin
				q			<=			16'hFFF0;
		end
		32'h00003304: begin
				q			<=			16'h16E3;
		end
		32'h00003306: begin
				q			<=			16'h66FB;
		end
		32'h00003308: begin
				q			<=			16'h98E3;
		end
		32'h0000330A: begin
				q			<=			16'h6E0C;
		end
		32'h0000330C: begin
				q			<=			16'h0793;
		end
		32'h0000330E: begin
				q			<=			16'h0090;
		end
		32'h00003310: begin
				q			<=			16'hE4E3;
		end
		32'h00003312: begin
				q			<=			16'h6F87;
		end
		32'h00003314: begin
				q			<=			16'h0C13;
		end
		32'h00003316: begin
				q			<=			16'h030C;
		end
		32'h00003318: begin
				q			<=			16'h07A3;
		end
		32'h0000331A: begin
				q			<=			16'h1981;
		end
		32'h0000331C: begin
				q			<=			16'h0493;
		end
		32'h0000331E: begin
				q			<=			16'h18F1;
		end
		32'h00003320: begin
				q			<=			16'h006F;
		end
		32'h00003322: begin
				q			<=			16'h6B10;
		end
		32'h00003324: begin
				q			<=			16'h8793;
		end
		32'h00003326: begin
				q			<=			16'h004A;
		end
		32'h00003328: begin
				q			<=			16'h2623;
		end
		32'h0000332A: begin
				q			<=			16'h00F1;
		end
		32'h0000332C: begin
				q			<=			16'h7793;
		end
		32'h0000332E: begin
				q			<=			16'h0104;
		end
		32'h00003330: begin
				q			<=			16'h8863;
		end
		32'h00003332: begin
				q			<=			16'h0007;
		end
		32'h00003334: begin
				q			<=			16'hAC03;
		end
		32'h00003336: begin
				q			<=			16'h000A;
		end
		32'h00003338: begin
				q			<=			16'h5C93;
		end
		32'h0000333A: begin
				q			<=			16'h41FC;
		end
		32'h0000333C: begin
				q			<=			16'hF06F;
		end
		32'h0000333E: begin
				q			<=			16'hFA9F;
		end
		32'h00003340: begin
				q			<=			16'h7793;
		end
		32'h00003342: begin
				q			<=			16'h0404;
		end
		32'h00003344: begin
				q			<=			16'hAC03;
		end
		32'h00003346: begin
				q			<=			16'h000A;
		end
		32'h00003348: begin
				q			<=			16'h8863;
		end
		32'h0000334A: begin
				q			<=			16'h0007;
		end
		32'h0000334C: begin
				q			<=			16'h1C13;
		end
		32'h0000334E: begin
				q			<=			16'h010C;
		end
		32'h00003350: begin
				q			<=			16'h5C13;
		end
		32'h00003352: begin
				q			<=			16'h410C;
		end
		32'h00003354: begin
				q			<=			16'hF06F;
		end
		32'h00003356: begin
				q			<=			16'hFE5F;
		end
		32'h00003358: begin
				q			<=			16'h7793;
		end
		32'h0000335A: begin
				q			<=			16'h2004;
		end
		32'h0000335C: begin
				q			<=			16'h8EE3;
		end
		32'h0000335E: begin
				q			<=			16'hFC07;
		end
		32'h00003360: begin
				q			<=			16'h1C13;
		end
		32'h00003362: begin
				q			<=			16'h018C;
		end
		32'h00003364: begin
				q			<=			16'h5C13;
		end
		32'h00003366: begin
				q			<=			16'h418C;
		end
		32'h00003368: begin
				q			<=			16'hF06F;
		end
		32'h0000336A: begin
				q			<=			16'hFD1F;
		end
		32'h0000336C: begin
				q			<=			16'h7793;
		end
		32'h0000336E: begin
				q			<=			16'h0084;
		end
		32'h00003370: begin
				q			<=			16'h8263;
		end
		32'h00003372: begin
				q			<=			16'h0C07;
		end
		32'h00003374: begin
				q			<=			16'h8793;
		end
		32'h00003376: begin
				q			<=			16'h004A;
		end
		32'h00003378: begin
				q			<=			16'h2623;
		end
		32'h0000337A: begin
				q			<=			16'h00F1;
		end
		32'h0000337C: begin
				q			<=			16'hA783;
		end
		32'h0000337E: begin
				q			<=			16'h000A;
		end
		32'h00003380: begin
				q			<=			16'hA603;
		end
		32'h00003382: begin
				q			<=			16'h0007;
		end
		32'h00003384: begin
				q			<=			16'hA683;
		end
		32'h00003386: begin
				q			<=			16'h0047;
		end
		32'h00003388: begin
				q			<=			16'hA703;
		end
		32'h0000338A: begin
				q			<=			16'h0087;
		end
		32'h0000338C: begin
				q			<=			16'hA783;
		end
		32'h0000338E: begin
				q			<=			16'h00C7;
		end
		32'h00003390: begin
				q			<=			16'h2823;
		end
		32'h00003392: begin
				q			<=			16'h0CC1;
		end
		32'h00003394: begin
				q			<=			16'h2A23;
		end
		32'h00003396: begin
				q			<=			16'h0CD1;
		end
		32'h00003398: begin
				q			<=			16'h2C23;
		end
		32'h0000339A: begin
				q			<=			16'h0CE1;
		end
		32'h0000339C: begin
				q			<=			16'h2E23;
		end
		32'h0000339E: begin
				q			<=			16'h0CF1;
		end
		32'h000033A0: begin
				q			<=			16'h0513;
		end
		32'h000033A2: begin
				q			<=			16'h0D01;
		end
		32'h000033A4: begin
				q			<=			16'h2223;
		end
		32'h000033A6: begin
				q			<=			16'h0111;
		end
		32'h000033A8: begin
				q			<=			16'h30EF;
		end
		32'h000033AA: begin
				q			<=			16'h73D0;
		end
		32'h000033AC: begin
				q			<=			16'h2623;
		end
		32'h000033AE: begin
				q			<=			16'h0AA1;
		end
		32'h000033B0: begin
				q			<=			16'h0793;
		end
		32'h000033B2: begin
				q			<=			16'h0020;
		end
		32'h000033B4: begin
				q			<=			16'h2883;
		end
		32'h000033B6: begin
				q			<=			16'h0041;
		end
		32'h000033B8: begin
				q			<=			16'h1463;
		end
		32'h000033BA: begin
				q			<=			16'h0CF5;
		end
		32'h000033BC: begin
				q			<=			16'h2783;
		end
		32'h000033BE: begin
				q			<=			16'h0D01;
		end
		32'h000033C0: begin
				q			<=			16'h0593;
		end
		32'h000033C2: begin
				q			<=			16'h0801;
		end
		32'h000033C4: begin
				q			<=			16'h0513;
		end
		32'h000033C6: begin
				q			<=			16'h0901;
		end
		32'h000033C8: begin
				q			<=			16'h2823;
		end
		32'h000033CA: begin
				q			<=			16'h08F1;
		end
		32'h000033CC: begin
				q			<=			16'h2783;
		end
		32'h000033CE: begin
				q			<=			16'h0D41;
		end
		32'h000033D0: begin
				q			<=			16'h2023;
		end
		32'h000033D2: begin
				q			<=			16'h0801;
		end
		32'h000033D4: begin
				q			<=			16'h2223;
		end
		32'h000033D6: begin
				q			<=			16'h0801;
		end
		32'h000033D8: begin
				q			<=			16'h2A23;
		end
		32'h000033DA: begin
				q			<=			16'h08F1;
		end
		32'h000033DC: begin
				q			<=			16'h2783;
		end
		32'h000033DE: begin
				q			<=			16'h0D81;
		end
		32'h000033E0: begin
				q			<=			16'h2423;
		end
		32'h000033E2: begin
				q			<=			16'h0801;
		end
		32'h000033E4: begin
				q			<=			16'h2623;
		end
		32'h000033E6: begin
				q			<=			16'h0801;
		end
		32'h000033E8: begin
				q			<=			16'h2C23;
		end
		32'h000033EA: begin
				q			<=			16'h08F1;
		end
		32'h000033EC: begin
				q			<=			16'h2783;
		end
		32'h000033EE: begin
				q			<=			16'h0DC1;
		end
		32'h000033F0: begin
				q			<=			16'h2E23;
		end
		32'h000033F2: begin
				q			<=			16'h08F1;
		end
		32'h000033F4: begin
				q			<=			16'h80EF;
		end
		32'h000033F6: begin
				q			<=			16'h5FD0;
		end
		32'h000033F8: begin
				q			<=			16'h2883;
		end
		32'h000033FA: begin
				q			<=			16'h0041;
		end
		32'h000033FC: begin
				q			<=			16'h5663;
		end
		32'h000033FE: begin
				q			<=			16'h0005;
		end
		32'h00003400: begin
				q			<=			16'h0793;
		end
		32'h00003402: begin
				q			<=			16'h02D0;
		end
		32'h00003404: begin
				q			<=			16'h03A3;
		end
		32'h00003406: begin
				q			<=			16'h0AF1;
		end
		32'h00003408: begin
				q			<=			16'h0793;
		end
		32'h0000340A: begin
				q			<=			16'h0470;
		end
		32'h0000340C: begin
				q			<=			16'hD497;
		end
		32'h0000340E: begin
				q			<=			16'h0000;
		end
		32'h00003410: begin
				q			<=			16'h8493;
		end
		32'h00003412: begin
				q			<=			16'h96C4;
		end
		32'h00003414: begin
				q			<=			16'hC663;
		end
		32'h00003416: begin
				q			<=			16'h01A7;
		end
		32'h00003418: begin
				q			<=			16'hD497;
		end
		32'h0000341A: begin
				q			<=			16'h0000;
		end
		32'h0000341C: begin
				q			<=			16'h8493;
		end
		32'h0000341E: begin
				q			<=			16'h95C4;
		end
		32'h00003420: begin
				q			<=			16'h7413;
		end
		32'h00003422: begin
				q			<=			16'hF7F4;
		end
		32'h00003424: begin
				q			<=			16'h2223;
		end
		32'h00003426: begin
				q			<=			16'h0001;
		end
		32'h00003428: begin
				q			<=			16'h0B13;
		end
		32'h0000342A: begin
				q			<=			16'h0030;
		end
		32'h0000342C: begin
				q			<=			16'h0D93;
		end
		32'h0000342E: begin
				q			<=			16'h0000;
		end
		32'h00003430: begin
				q			<=			16'h006F;
		end
		32'h00003432: begin
				q			<=			16'h5B10;
		end
		32'h00003434: begin
				q			<=			16'h8A93;
		end
		32'h00003436: begin
				q			<=			16'h007A;
		end
		32'h00003438: begin
				q			<=			16'hFA93;
		end
		32'h0000343A: begin
				q			<=			16'hFF8A;
		end
		32'h0000343C: begin
				q			<=			16'hA583;
		end
		32'h0000343E: begin
				q			<=			16'h000A;
		end
		32'h00003440: begin
				q			<=			16'hA603;
		end
		32'h00003442: begin
				q			<=			16'h004A;
		end
		32'h00003444: begin
				q			<=			16'h8793;
		end
		32'h00003446: begin
				q			<=			16'h008A;
		end
		32'h00003448: begin
				q			<=			16'h0513;
		end
		32'h0000344A: begin
				q			<=			16'h0901;
		end
		32'h0000344C: begin
				q			<=			16'h2223;
		end
		32'h0000344E: begin
				q			<=			16'h0111;
		end
		32'h00003450: begin
				q			<=			16'h2623;
		end
		32'h00003452: begin
				q			<=			16'h00F1;
		end
		32'h00003454: begin
				q			<=			16'hB0EF;
		end
		32'h00003456: begin
				q			<=			16'h6F40;
		end
		32'h00003458: begin
				q			<=			16'h2783;
		end
		32'h0000345A: begin
				q			<=			16'h0901;
		end
		32'h0000345C: begin
				q			<=			16'h2883;
		end
		32'h0000345E: begin
				q			<=			16'h0041;
		end
		32'h00003460: begin
				q			<=			16'h2823;
		end
		32'h00003462: begin
				q			<=			16'h0CF1;
		end
		32'h00003464: begin
				q			<=			16'h2783;
		end
		32'h00003466: begin
				q			<=			16'h0941;
		end
		32'h00003468: begin
				q			<=			16'h2A23;
		end
		32'h0000346A: begin
				q			<=			16'h0CF1;
		end
		32'h0000346C: begin
				q			<=			16'h2783;
		end
		32'h0000346E: begin
				q			<=			16'h0981;
		end
		32'h00003470: begin
				q			<=			16'h2C23;
		end
		32'h00003472: begin
				q			<=			16'h0CF1;
		end
		32'h00003474: begin
				q			<=			16'h2783;
		end
		32'h00003476: begin
				q			<=			16'h09C1;
		end
		32'h00003478: begin
				q			<=			16'h2E23;
		end
		32'h0000347A: begin
				q			<=			16'h0CF1;
		end
		32'h0000347C: begin
				q			<=			16'hF06F;
		end
		32'h0000347E: begin
				q			<=			16'hF25F;
		end
		32'h00003480: begin
				q			<=			16'h0793;
		end
		32'h00003482: begin
				q			<=			16'h0010;
		end
		32'h00003484: begin
				q			<=			16'h1063;
		end
		32'h00003486: begin
				q			<=			16'h02F5;
		end
		32'h00003488: begin
				q			<=			16'h0793;
		end
		32'h0000348A: begin
				q			<=			16'h0470;
		end
		32'h0000348C: begin
				q			<=			16'hD497;
		end
		32'h0000348E: begin
				q			<=			16'h0000;
		end
		32'h00003490: begin
				q			<=			16'h8493;
		end
		32'h00003492: begin
				q			<=			16'h8F44;
		end
		32'h00003494: begin
				q			<=			16'hC6E3;
		end
		32'h00003496: begin
				q			<=			16'hF9A7;
		end
		32'h00003498: begin
				q			<=			16'hD497;
		end
		32'h0000349A: begin
				q			<=			16'h0000;
		end
		32'h0000349C: begin
				q			<=			16'h8493;
		end
		32'h0000349E: begin
				q			<=			16'h8E44;
		end
		32'h000034A0: begin
				q			<=			16'hF06F;
		end
		32'h000034A2: begin
				q			<=			16'hF81F;
		end
		32'h000034A4: begin
				q			<=			16'h7B93;
		end
		32'h000034A6: begin
				q			<=			16'hFDFD;
		end
		32'h000034A8: begin
				q			<=			16'h0793;
		end
		32'h000034AA: begin
				q			<=			16'h0410;
		end
		32'h000034AC: begin
				q			<=			16'h9063;
		end
		32'h000034AE: begin
				q			<=			16'h0AFB;
		end
		32'h000034B0: begin
				q			<=			16'h0793;
		end
		32'h000034B2: begin
				q			<=			16'h0300;
		end
		32'h000034B4: begin
				q			<=			16'h0423;
		end
		32'h000034B6: begin
				q			<=			16'h0AF1;
		end
		32'h000034B8: begin
				q			<=			16'h0713;
		end
		32'h000034BA: begin
				q			<=			16'h0610;
		end
		32'h000034BC: begin
				q			<=			16'h0793;
		end
		32'h000034BE: begin
				q			<=			16'h0580;
		end
		32'h000034C0: begin
				q			<=			16'h1463;
		end
		32'h000034C2: begin
				q			<=			16'h00ED;
		end
		32'h000034C4: begin
				q			<=			16'h0793;
		end
		32'h000034C6: begin
				q			<=			16'h0780;
		end
		32'h000034C8: begin
				q			<=			16'h04A3;
		end
		32'h000034CA: begin
				q			<=			16'h0AF1;
		end
		32'h000034CC: begin
				q			<=			16'h0793;
		end
		32'h000034CE: begin
				q			<=			16'h0630;
		end
		32'h000034D0: begin
				q			<=			16'h6413;
		end
		32'h000034D2: begin
				q			<=			16'h0024;
		end
		32'h000034D4: begin
				q			<=			16'hD663;
		end
		32'h000034D6: begin
				q			<=			16'h4F67;
		end
		32'h000034D8: begin
				q			<=			16'h0593;
		end
		32'h000034DA: begin
				q			<=			16'h001B;
		end
		32'h000034DC: begin
				q			<=			16'h0513;
		end
		32'h000034DE: begin
				q			<=			16'h0009;
		end
		32'h000034E0: begin
				q			<=			16'h2223;
		end
		32'h000034E2: begin
				q			<=			16'h0111;
		end
		32'h000034E4: begin
				q			<=			16'h30EF;
		end
		32'h000034E6: begin
				q			<=			16'h6BD0;
		end
		32'h000034E8: begin
				q			<=			16'h0493;
		end
		32'h000034EA: begin
				q			<=			16'h0005;
		end
		32'h000034EC: begin
				q			<=			16'h2883;
		end
		32'h000034EE: begin
				q			<=			16'h0041;
		end
		32'h000034F0: begin
				q			<=			16'h1E63;
		end
		32'h000034F2: begin
				q			<=			16'h4C05;
		end
		32'h000034F4: begin
				q			<=			16'hD783;
		end
		32'h000034F6: begin
				q			<=			16'h00C9;
		end
		32'h000034F8: begin
				q			<=			16'hE793;
		end
		32'h000034FA: begin
				q			<=			16'h0407;
		end
		32'h000034FC: begin
				q			<=			16'h9623;
		end
		32'h000034FE: begin
				q			<=			16'h00F9;
		end
		32'h00003500: begin
				q			<=			16'hD783;
		end
		32'h00003502: begin
				q			<=			16'h00C9;
		end
		32'h00003504: begin
				q			<=			16'hF793;
		end
		32'h00003506: begin
				q			<=			16'h0407;
		end
		32'h00003508: begin
				q			<=			16'h9CE3;
		end
		32'h0000350A: begin
				q			<=			16'hA607;
		end
		32'h0000350C: begin
				q			<=			16'h2083;
		end
		32'h0000350E: begin
				q			<=			16'h1CC1;
		end
		32'h00003510: begin
				q			<=			16'h2403;
		end
		32'h00003512: begin
				q			<=			16'h1C81;
		end
		32'h00003514: begin
				q			<=			16'h2503;
		end
		32'h00003516: begin
				q			<=			16'h0181;
		end
		32'h00003518: begin
				q			<=			16'h2483;
		end
		32'h0000351A: begin
				q			<=			16'h1C41;
		end
		32'h0000351C: begin
				q			<=			16'h2903;
		end
		32'h0000351E: begin
				q			<=			16'h1C01;
		end
		32'h00003520: begin
				q			<=			16'h2983;
		end
		32'h00003522: begin
				q			<=			16'h1BC1;
		end
		32'h00003524: begin
				q			<=			16'h2A03;
		end
		32'h00003526: begin
				q			<=			16'h1B81;
		end
		32'h00003528: begin
				q			<=			16'h2A83;
		end
		32'h0000352A: begin
				q			<=			16'h1B41;
		end
		32'h0000352C: begin
				q			<=			16'h2B03;
		end
		32'h0000352E: begin
				q			<=			16'h1B01;
		end
		32'h00003530: begin
				q			<=			16'h2B83;
		end
		32'h00003532: begin
				q			<=			16'h1AC1;
		end
		32'h00003534: begin
				q			<=			16'h2C03;
		end
		32'h00003536: begin
				q			<=			16'h1A81;
		end
		32'h00003538: begin
				q			<=			16'h2C83;
		end
		32'h0000353A: begin
				q			<=			16'h1A41;
		end
		32'h0000353C: begin
				q			<=			16'h2D03;
		end
		32'h0000353E: begin
				q			<=			16'h1A01;
		end
		32'h00003540: begin
				q			<=			16'h2D83;
		end
		32'h00003542: begin
				q			<=			16'h19C1;
		end
		32'h00003544: begin
				q			<=			16'h0113;
		end
		32'h00003546: begin
				q			<=			16'h1D01;
		end
		32'h00003548: begin
				q			<=			16'h8067;
		end
		32'h0000354A: begin
				q			<=			16'h0000;
		end
		32'h0000354C: begin
				q			<=			16'h0793;
		end
		32'h0000354E: begin
				q			<=			16'hFFF0;
		end
		32'h00003550: begin
				q			<=			16'h0263;
		end
		32'h00003552: begin
				q			<=			16'h48FB;
		end
		32'h00003554: begin
				q			<=			16'h0793;
		end
		32'h00003556: begin
				q			<=			16'h0470;
		end
		32'h00003558: begin
				q			<=			16'h2223;
		end
		32'h0000355A: begin
				q			<=			16'h0001;
		end
		32'h0000355C: begin
				q			<=			16'h9463;
		end
		32'h0000355E: begin
				q			<=			16'h00FB;
		end
		32'h00003560: begin
				q			<=			16'h0063;
		end
		32'h00003562: begin
				q			<=			16'h480B;
		end
		32'h00003564: begin
				q			<=			16'h2A83;
		end
		32'h00003566: begin
				q			<=			16'h0DC1;
		end
		32'h00003568: begin
				q			<=			16'h6793;
		end
		32'h0000356A: begin
				q			<=			16'h1004;
		end
		32'h0000356C: begin
				q			<=			16'h2023;
		end
		32'h0000356E: begin
				q			<=			16'h02F1;
		end
		32'h00003570: begin
				q			<=			16'h2C23;
		end
		32'h00003572: begin
				q			<=			16'h0201;
		end
		32'h00003574: begin
				q			<=			16'h2E03;
		end
		32'h00003576: begin
				q			<=			16'h0D01;
		end
		32'h00003578: begin
				q			<=			16'h2D83;
		end
		32'h0000357A: begin
				q			<=			16'h0D41;
		end
		32'h0000357C: begin
				q			<=			16'h2C83;
		end
		32'h0000357E: begin
				q			<=			16'h0D81;
		end
		32'h00003580: begin
				q			<=			16'hDA63;
		end
		32'h00003582: begin
				q			<=			16'h000A;
		end
		32'h00003584: begin
				q			<=			16'h07B7;
		end
		32'h00003586: begin
				q			<=			16'h8000;
		end
		32'h00003588: begin
				q			<=			16'hCAB3;
		end
		32'h0000358A: begin
				q			<=			16'h0157;
		end
		32'h0000358C: begin
				q			<=			16'h0793;
		end
		32'h0000358E: begin
				q			<=			16'h02D0;
		end
		32'h00003590: begin
				q			<=			16'h2C23;
		end
		32'h00003592: begin
				q			<=			16'h02F1;
		end
		32'h00003594: begin
				q			<=			16'h0793;
		end
		32'h00003596: begin
				q			<=			16'h0410;
		end
		32'h00003598: begin
				q			<=			16'h9863;
		end
		32'h0000359A: begin
				q			<=			16'h48FB;
		end
		32'h0000359C: begin
				q			<=			16'h0513;
		end
		32'h0000359E: begin
				q			<=			16'h0901;
		end
		32'h000035A0: begin
				q			<=			16'h2423;
		end
		32'h000035A2: begin
				q			<=			16'h0511;
		end
		32'h000035A4: begin
				q			<=			16'h2823;
		end
		32'h000035A6: begin
				q			<=			16'h09C1;
		end
		32'h000035A8: begin
				q			<=			16'h2C23;
		end
		32'h000035AA: begin
				q			<=			16'h0991;
		end
		32'h000035AC: begin
				q			<=			16'h2A23;
		end
		32'h000035AE: begin
				q			<=			16'h09B1;
		end
		32'h000035B0: begin
				q			<=			16'h2E23;
		end
		32'h000035B2: begin
				q			<=			16'h0951;
		end
		32'h000035B4: begin
				q			<=			16'hB0EF;
		end
		32'h000035B6: begin
				q			<=			16'h7BC0;
		end
		32'h000035B8: begin
				q			<=			16'h0613;
		end
		32'h000035BA: begin
				q			<=			16'h0AC1;
		end
		32'h000035BC: begin
				q			<=			16'h50EF;
		end
		32'h000035BE: begin
				q			<=			16'h3940;
		end
		32'h000035C0: begin
				q			<=			16'h8613;
		end
		32'h000035C2: begin
				q			<=			16'h0005;
		end
		32'h000035C4: begin
				q			<=			16'h0593;
		end
		32'h000035C6: begin
				q			<=			16'h0005;
		end
		32'h000035C8: begin
				q			<=			16'h0513;
		end
		32'h000035CA: begin
				q			<=			16'h0901;
		end
		32'h000035CC: begin
				q			<=			16'hB0EF;
		end
		32'h000035CE: begin
				q			<=			16'h57C0;
		end
		32'h000035D0: begin
				q			<=			16'h2783;
		end
		32'h000035D2: begin
				q			<=			16'h0901;
		end
		32'h000035D4: begin
				q			<=			16'h0613;
		end
		32'h000035D6: begin
				q			<=			16'h0601;
		end
		32'h000035D8: begin
				q			<=			16'h0593;
		end
		32'h000035DA: begin
				q			<=			16'h0701;
		end
		32'h000035DC: begin
				q			<=			16'h2823;
		end
		32'h000035DE: begin
				q			<=			16'h06F1;
		end
		32'h000035E0: begin
				q			<=			16'h2783;
		end
		32'h000035E2: begin
				q			<=			16'h0941;
		end
		32'h000035E4: begin
				q			<=			16'h0513;
		end
		32'h000035E6: begin
				q			<=			16'h0801;
		end
		32'h000035E8: begin
				q			<=			16'h2023;
		end
		32'h000035EA: begin
				q			<=			16'h0601;
		end
		32'h000035EC: begin
				q			<=			16'h2A23;
		end
		32'h000035EE: begin
				q			<=			16'h06F1;
		end
		32'h000035F0: begin
				q			<=			16'h2783;
		end
		32'h000035F2: begin
				q			<=			16'h0981;
		end
		32'h000035F4: begin
				q			<=			16'h2223;
		end
		32'h000035F6: begin
				q			<=			16'h0601;
		end
		32'h000035F8: begin
				q			<=			16'h2423;
		end
		32'h000035FA: begin
				q			<=			16'h0601;
		end
		32'h000035FC: begin
				q			<=			16'h2C23;
		end
		32'h000035FE: begin
				q			<=			16'h06F1;
		end
		32'h00003600: begin
				q			<=			16'h2783;
		end
		32'h00003602: begin
				q			<=			16'h09C1;
		end
		32'h00003604: begin
				q			<=			16'h2E23;
		end
		32'h00003606: begin
				q			<=			16'h06F1;
		end
		32'h00003608: begin
				q			<=			16'h07B7;
		end
		32'h0000360A: begin
				q			<=			16'h3FFC;
		end
		32'h0000360C: begin
				q			<=			16'h2623;
		end
		32'h0000360E: begin
				q			<=			16'h06F1;
		end
		32'h00003610: begin
				q			<=			16'h80EF;
		end
		32'h00003612: begin
				q			<=			16'h5450;
		end
		32'h00003614: begin
				q			<=			16'h2803;
		end
		32'h00003616: begin
				q			<=			16'h0801;
		end
		32'h00003618: begin
				q			<=			16'h2603;
		end
		32'h0000361A: begin
				q			<=			16'h0841;
		end
		32'h0000361C: begin
				q			<=			16'h2683;
		end
		32'h0000361E: begin
				q			<=			16'h0881;
		end
		32'h00003620: begin
				q			<=			16'h2C83;
		end
		32'h00003622: begin
				q			<=			16'h08C1;
		end
		32'h00003624: begin
				q			<=			16'h0593;
		end
		32'h00003626: begin
				q			<=			16'h0801;
		end
		32'h00003628: begin
				q			<=			16'h0513;
		end
		32'h0000362A: begin
				q			<=			16'h0901;
		end
		32'h0000362C: begin
				q			<=			16'h2823;
		end
		32'h0000362E: begin
				q			<=			16'h0901;
		end
		32'h00003630: begin
				q			<=			16'h2223;
		end
		32'h00003632: begin
				q			<=			16'h0501;
		end
		32'h00003634: begin
				q			<=			16'h2A23;
		end
		32'h00003636: begin
				q			<=			16'h08C1;
		end
		32'h00003638: begin
				q			<=			16'h2023;
		end
		32'h0000363A: begin
				q			<=			16'h04C1;
		end
		32'h0000363C: begin
				q			<=			16'h2C23;
		end
		32'h0000363E: begin
				q			<=			16'h08D1;
		end
		32'h00003640: begin
				q			<=			16'h2E23;
		end
		32'h00003642: begin
				q			<=			16'h02D1;
		end
		32'h00003644: begin
				q			<=			16'h2E23;
		end
		32'h00003646: begin
				q			<=			16'h0991;
		end
		32'h00003648: begin
				q			<=			16'h2023;
		end
		32'h0000364A: begin
				q			<=			16'h0801;
		end
		32'h0000364C: begin
				q			<=			16'h2223;
		end
		32'h0000364E: begin
				q			<=			16'h0801;
		end
		32'h00003650: begin
				q			<=			16'h2423;
		end
		32'h00003652: begin
				q			<=			16'h0801;
		end
		32'h00003654: begin
				q			<=			16'h2623;
		end
		32'h00003656: begin
				q			<=			16'h0801;
		end
		32'h00003658: begin
				q			<=			16'h80EF;
		end
		32'h0000365A: begin
				q			<=			16'h1650;
		end
		32'h0000365C: begin
				q			<=			16'h2683;
		end
		32'h0000365E: begin
				q			<=			16'h03C1;
		end
		32'h00003660: begin
				q			<=			16'h2603;
		end
		32'h00003662: begin
				q			<=			16'h0401;
		end
		32'h00003664: begin
				q			<=			16'h2803;
		end
		32'h00003666: begin
				q			<=			16'h0441;
		end
		32'h00003668: begin
				q			<=			16'h2883;
		end
		32'h0000366A: begin
				q			<=			16'h0481;
		end
		32'h0000366C: begin
				q			<=			16'h1663;
		end
		32'h0000366E: begin
				q			<=			16'h0005;
		end
		32'h00003670: begin
				q			<=			16'h0713;
		end
		32'h00003672: begin
				q			<=			16'h0010;
		end
		32'h00003674: begin
				q			<=			16'h2623;
		end
		32'h00003676: begin
				q			<=			16'h0AE1;
		end
		32'h00003678: begin
				q			<=			16'h0713;
		end
		32'h0000367A: begin
				q			<=			16'h0610;
		end
		32'h0000367C: begin
				q			<=			16'hCA97;
		end
		32'h0000367E: begin
				q			<=			16'h0000;
		end
		32'h00003680: begin
				q			<=			16'h8A93;
		end
		32'h00003682: begin
				q			<=			16'h71CA;
		end
		32'h00003684: begin
				q			<=			16'h1663;
		end
		32'h00003686: begin
				q			<=			16'h00ED;
		end
		32'h00003688: begin
				q			<=			16'hCA97;
		end
		32'h0000368A: begin
				q			<=			16'h0000;
		end
		32'h0000368C: begin
				q			<=			16'h8A93;
		end
		32'h0000368E: begin
				q			<=			16'h6FCA;
		end
		32'h00003690: begin
				q			<=			16'h0E13;
		end
		32'h00003692: begin
				q			<=			16'hFFFB;
		end
		32'h00003694: begin
				q			<=			16'h8D93;
		end
		32'h00003696: begin
				q			<=			16'h0004;
		end
		32'h00003698: begin
				q			<=			16'h07B7;
		end
		32'h0000369A: begin
				q			<=			16'h4003;
		end
		32'h0000369C: begin
				q			<=			16'h0593;
		end
		32'h0000369E: begin
				q			<=			16'h0801;
		end
		32'h000036A0: begin
				q			<=			16'h2223;
		end
		32'h000036A2: begin
				q			<=			16'h08C1;
		end
		32'h000036A4: begin
				q			<=			16'h0513;
		end
		32'h000036A6: begin
				q			<=			16'h0901;
		end
		32'h000036A8: begin
				q			<=			16'h0613;
		end
		32'h000036AA: begin
				q			<=			16'h0701;
		end
		32'h000036AC: begin
				q			<=			16'h2423;
		end
		32'h000036AE: begin
				q			<=			16'h0511;
		end
		32'h000036B0: begin
				q			<=			16'h2223;
		end
		32'h000036B2: begin
				q			<=			16'h05C1;
		end
		32'h000036B4: begin
				q			<=			16'h2023;
		end
		32'h000036B6: begin
				q			<=			16'h0901;
		end
		32'h000036B8: begin
				q			<=			16'h2E23;
		end
		32'h000036BA: begin
				q			<=			16'h06F1;
		end
		32'h000036BC: begin
				q			<=			16'h2423;
		end
		32'h000036BE: begin
				q			<=			16'h08D1;
		end
		32'h000036C0: begin
				q			<=			16'h2623;
		end
		32'h000036C2: begin
				q			<=			16'h0991;
		end
		32'h000036C4: begin
				q			<=			16'h2823;
		end
		32'h000036C6: begin
				q			<=			16'h0601;
		end
		32'h000036C8: begin
				q			<=			16'h2A23;
		end
		32'h000036CA: begin
				q			<=			16'h0601;
		end
		32'h000036CC: begin
				q			<=			16'h2C23;
		end
		32'h000036CE: begin
				q			<=			16'h0601;
		end
		32'h000036D0: begin
				q			<=			16'h80EF;
		end
		32'h000036D2: begin
				q			<=			16'h4850;
		end
		32'h000036D4: begin
				q			<=			16'h2603;
		end
		32'h000036D6: begin
				q			<=			16'h0901;
		end
		32'h000036D8: begin
				q			<=			16'h2683;
		end
		32'h000036DA: begin
				q			<=			16'h0941;
		end
		32'h000036DC: begin
				q			<=			16'h0513;
		end
		32'h000036DE: begin
				q			<=			16'h0901;
		end
		32'h000036E0: begin
				q			<=			16'h2023;
		end
		32'h000036E2: begin
				q			<=			16'h04C1;
		end
		32'h000036E4: begin
				q			<=			16'h2E23;
		end
		32'h000036E6: begin
				q			<=			16'h02D1;
		end
		32'h000036E8: begin
				q			<=			16'hB0EF;
		end
		32'h000036EA: begin
				q			<=			16'h1740;
		end
		32'h000036EC: begin
				q			<=			16'h0593;
		end
		32'h000036EE: begin
				q			<=			16'h0005;
		end
		32'h000036F0: begin
				q			<=			16'h0A13;
		end
		32'h000036F2: begin
				q			<=			16'h0005;
		end
		32'h000036F4: begin
				q			<=			16'h0513;
		end
		32'h000036F6: begin
				q			<=			16'h0901;
		end
		32'h000036F8: begin
				q			<=			16'h2C83;
		end
		32'h000036FA: begin
				q			<=			16'h0981;
		end
		32'h000036FC: begin
				q			<=			16'h2C03;
		end
		32'h000036FE: begin
				q			<=			16'h09C1;
		end
		32'h00003700: begin
				q			<=			16'hB0EF;
		end
		32'h00003702: begin
				q			<=			16'h2C40;
		end
		32'h00003704: begin
				q			<=			16'h2783;
		end
		32'h00003706: begin
				q			<=			16'h0901;
		end
		32'h00003708: begin
				q			<=			16'h2603;
		end
		32'h0000370A: begin
				q			<=			16'h0401;
		end
		32'h0000370C: begin
				q			<=			16'h2683;
		end
		32'h0000370E: begin
				q			<=			16'h03C1;
		end
		32'h00003710: begin
				q			<=			16'h2023;
		end
		32'h00003712: begin
				q			<=			16'h06F1;
		end
		32'h00003714: begin
				q			<=			16'h2783;
		end
		32'h00003716: begin
				q			<=			16'h0941;
		end
		32'h00003718: begin
				q			<=			16'h2823;
		end
		32'h0000371A: begin
				q			<=			16'h06C1;
		end
		32'h0000371C: begin
				q			<=			16'h0593;
		end
		32'h0000371E: begin
				q			<=			16'h0701;
		end
		32'h00003720: begin
				q			<=			16'h2223;
		end
		32'h00003722: begin
				q			<=			16'h06F1;
		end
		32'h00003724: begin
				q			<=			16'h2783;
		end
		32'h00003726: begin
				q			<=			16'h0981;
		end
		32'h00003728: begin
				q			<=			16'h0613;
		end
		32'h0000372A: begin
				q			<=			16'h0601;
		end
		32'h0000372C: begin
				q			<=			16'h0513;
		end
		32'h0000372E: begin
				q			<=			16'h0801;
		end
		32'h00003730: begin
				q			<=			16'h2423;
		end
		32'h00003732: begin
				q			<=			16'h06F1;
		end
		32'h00003734: begin
				q			<=			16'h2783;
		end
		32'h00003736: begin
				q			<=			16'h09C1;
		end
		32'h00003738: begin
				q			<=			16'h2C23;
		end
		32'h0000373A: begin
				q			<=			16'h0791;
		end
		32'h0000373C: begin
				q			<=			16'h2E23;
		end
		32'h0000373E: begin
				q			<=			16'h0781;
		end
		32'h00003740: begin
				q			<=			16'h2623;
		end
		32'h00003742: begin
				q			<=			16'h06F1;
		end
		32'h00003744: begin
				q			<=			16'h2A23;
		end
		32'h00003746: begin
				q			<=			16'h06D1;
		end
		32'h00003748: begin
				q			<=			16'h90EF;
		end
		32'h0000374A: begin
				q			<=			16'h4510;
		end
		32'h0000374C: begin
				q			<=			16'h85B3;
		end
		32'h0000374E: begin
				q			<=			16'h014A;
		end
		32'h00003750: begin
				q			<=			16'hC583;
		end
		32'h00003752: begin
				q			<=			16'h0005;
		end
		32'h00003754: begin
				q			<=			16'h2E03;
		end
		32'h00003756: begin
				q			<=			16'h0441;
		end
		32'h00003758: begin
				q			<=			16'h2C03;
		end
		32'h0000375A: begin
				q			<=			16'h08C1;
		end
		32'h0000375C: begin
				q			<=			16'h8D93;
		end
		32'h0000375E: begin
				q			<=			16'h001D;
		end
		32'h00003760: begin
				q			<=			16'h2283;
		end
		32'h00003762: begin
				q			<=			16'h0801;
		end
		32'h00003764: begin
				q			<=			16'h2F83;
		end
		32'h00003766: begin
				q			<=			16'h0841;
		end
		32'h00003768: begin
				q			<=			16'h2F03;
		end
		32'h0000376A: begin
				q			<=			16'h0881;
		end
		32'h0000376C: begin
				q			<=			16'h2E23;
		end
		32'h0000376E: begin
				q			<=			16'h03C1;
		end
		32'h00003770: begin
				q			<=			16'h8FA3;
		end
		32'h00003772: begin
				q			<=			16'hFEBD;
		end
		32'h00003774: begin
				q			<=			16'h0793;
		end
		32'h00003776: begin
				q			<=			16'hFFF0;
		end
		32'h00003778: begin
				q			<=			16'h0C93;
		end
		32'h0000377A: begin
				q			<=			16'h000C;
		end
		32'h0000377C: begin
				q			<=			16'h2883;
		end
		32'h0000377E: begin
				q			<=			16'h0481;
		end
		32'h00003780: begin
				q			<=			16'h0C63;
		end
		32'h00003782: begin
				q			<=			16'h06FE;
		end
		32'h00003784: begin
				q			<=			16'h0E13;
		end
		32'h00003786: begin
				q			<=			16'hFFFE;
		end
		32'h00003788: begin
				q			<=			16'h0593;
		end
		32'h0000378A: begin
				q			<=			16'h0801;
		end
		32'h0000378C: begin
				q			<=			16'h0513;
		end
		32'h0000378E: begin
				q			<=			16'h0901;
		end
		32'h00003790: begin
				q			<=			16'h2E23;
		end
		32'h00003792: begin
				q			<=			16'h05E1;
		end
		32'h00003794: begin
				q			<=			16'h2C23;
		end
		32'h00003796: begin
				q			<=			16'h05F1;
		end
		32'h00003798: begin
				q			<=			16'h2A23;
		end
		32'h0000379A: begin
				q			<=			16'h0451;
		end
		32'h0000379C: begin
				q			<=			16'h2823;
		end
		32'h0000379E: begin
				q			<=			16'h0511;
		end
		32'h000037A0: begin
				q			<=			16'h2623;
		end
		32'h000037A2: begin
				q			<=			16'h05C1;
		end
		32'h000037A4: begin
				q			<=			16'h2823;
		end
		32'h000037A6: begin
				q			<=			16'h0851;
		end
		32'h000037A8: begin
				q			<=			16'h2423;
		end
		32'h000037AA: begin
				q			<=			16'h0451;
		end
		32'h000037AC: begin
				q			<=			16'h2A23;
		end
		32'h000037AE: begin
				q			<=			16'h09F1;
		end
		32'h000037B0: begin
				q			<=			16'h2223;
		end
		32'h000037B2: begin
				q			<=			16'h05F1;
		end
		32'h000037B4: begin
				q			<=			16'h2C23;
		end
		32'h000037B6: begin
				q			<=			16'h09E1;
		end
		32'h000037B8: begin
				q			<=			16'h2023;
		end
		32'h000037BA: begin
				q			<=			16'h05E1;
		end
		32'h000037BC: begin
				q			<=			16'h2E23;
		end
		32'h000037BE: begin
				q			<=			16'h0981;
		end
		32'h000037C0: begin
				q			<=			16'h2023;
		end
		32'h000037C2: begin
				q			<=			16'h0801;
		end
		32'h000037C4: begin
				q			<=			16'h2223;
		end
		32'h000037C6: begin
				q			<=			16'h0801;
		end
		32'h000037C8: begin
				q			<=			16'h2423;
		end
		32'h000037CA: begin
				q			<=			16'h0801;
		end
		32'h000037CC: begin
				q			<=			16'h2623;
		end
		32'h000037CE: begin
				q			<=			16'h0801;
		end
		32'h000037D0: begin
				q			<=			16'h80EF;
		end
		32'h000037D2: begin
				q			<=			16'h7EC0;
		end
		32'h000037D4: begin
				q			<=			16'h2683;
		end
		32'h000037D6: begin
				q			<=			16'h0401;
		end
		32'h000037D8: begin
				q			<=			16'h2603;
		end
		32'h000037DA: begin
				q			<=			16'h0441;
		end
		32'h000037DC: begin
				q			<=			16'h2803;
		end
		32'h000037DE: begin
				q			<=			16'h0481;
		end
		32'h000037E0: begin
				q			<=			16'h2E03;
		end
		32'h000037E2: begin
				q			<=			16'h04C1;
		end
		32'h000037E4: begin
				q			<=			16'h2883;
		end
		32'h000037E6: begin
				q			<=			16'h0501;
		end
		32'h000037E8: begin
				q			<=			16'h2283;
		end
		32'h000037EA: begin
				q			<=			16'h0541;
		end
		32'h000037EC: begin
				q			<=			16'h2F83;
		end
		32'h000037EE: begin
				q			<=			16'h0581;
		end
		32'h000037F0: begin
				q			<=			16'h2F03;
		end
		32'h000037F2: begin
				q			<=			16'h05C1;
		end
		32'h000037F4: begin
				q			<=			16'h12E3;
		end
		32'h000037F6: begin
				q			<=			16'hEA05;
		end
		32'h000037F8: begin
				q			<=			16'h0CB7;
		end
		32'h000037FA: begin
				q			<=			16'h3FFE;
		end
		32'h000037FC: begin
				q			<=			16'h0593;
		end
		32'h000037FE: begin
				q			<=			16'h0801;
		end
		32'h00003800: begin
				q			<=			16'h0513;
		end
		32'h00003802: begin
				q			<=			16'h0901;
		end
		32'h00003804: begin
				q			<=			16'h2023;
		end
		32'h00003806: begin
				q			<=			16'h0511;
		end
		32'h00003808: begin
				q			<=			16'h2823;
		end
		32'h0000380A: begin
				q			<=			16'h0851;
		end
		32'h0000380C: begin
				q			<=			16'h2623;
		end
		32'h0000380E: begin
				q			<=			16'h0451;
		end
		32'h00003810: begin
				q			<=			16'h2A23;
		end
		32'h00003812: begin
				q			<=			16'h09F1;
		end
		32'h00003814: begin
				q			<=			16'h2423;
		end
		32'h00003816: begin
				q			<=			16'h05F1;
		end
		32'h00003818: begin
				q			<=			16'h2C23;
		end
		32'h0000381A: begin
				q			<=			16'h09E1;
		end
		32'h0000381C: begin
				q			<=			16'h2223;
		end
		32'h0000381E: begin
				q			<=			16'h05E1;
		end
		32'h00003820: begin
				q			<=			16'h2E23;
		end
		32'h00003822: begin
				q			<=			16'h0981;
		end
		32'h00003824: begin
				q			<=			16'h2023;
		end
		32'h00003826: begin
				q			<=			16'h0801;
		end
		32'h00003828: begin
				q			<=			16'h2223;
		end
		32'h0000382A: begin
				q			<=			16'h0801;
		end
		32'h0000382C: begin
				q			<=			16'h2423;
		end
		32'h0000382E: begin
				q			<=			16'h0801;
		end
		32'h00003830: begin
				q			<=			16'h2623;
		end
		32'h00003832: begin
				q			<=			16'h0991;
		end
		32'h00003834: begin
				q			<=			16'h80EF;
		end
		32'h00003836: begin
				q			<=			16'h0590;
		end
		32'h00003838: begin
				q			<=			16'h2883;
		end
		32'h0000383A: begin
				q			<=			16'h0401;
		end
		32'h0000383C: begin
				q			<=			16'h4663;
		end
		32'h0000383E: begin
				q			<=			16'h04A0;
		end
		32'h00003840: begin
				q			<=			16'h2283;
		end
		32'h00003842: begin
				q			<=			16'h04C1;
		end
		32'h00003844: begin
				q			<=			16'h2F83;
		end
		32'h00003846: begin
				q			<=			16'h0481;
		end
		32'h00003848: begin
				q			<=			16'h2F03;
		end
		32'h0000384A: begin
				q			<=			16'h0441;
		end
		32'h0000384C: begin
				q			<=			16'h0593;
		end
		32'h0000384E: begin
				q			<=			16'h0801;
		end
		32'h00003850: begin
				q			<=			16'h0513;
		end
		32'h00003852: begin
				q			<=			16'h0901;
		end
		32'h00003854: begin
				q			<=			16'h2823;
		end
		32'h00003856: begin
				q			<=			16'h0851;
		end
		32'h00003858: begin
				q			<=			16'h2A23;
		end
		32'h0000385A: begin
				q			<=			16'h09F1;
		end
		32'h0000385C: begin
				q			<=			16'h2C23;
		end
		32'h0000385E: begin
				q			<=			16'h09E1;
		end
		32'h00003860: begin
				q			<=			16'h2E23;
		end
		32'h00003862: begin
				q			<=			16'h0981;
		end
		32'h00003864: begin
				q			<=			16'h2023;
		end
		32'h00003866: begin
				q			<=			16'h0801;
		end
		32'h00003868: begin
				q			<=			16'h2223;
		end
		32'h0000386A: begin
				q			<=			16'h0801;
		end
		32'h0000386C: begin
				q			<=			16'h2423;
		end
		32'h0000386E: begin
				q			<=			16'h0801;
		end
		32'h00003870: begin
				q			<=			16'h2623;
		end
		32'h00003872: begin
				q			<=			16'h0991;
		end
		32'h00003874: begin
				q			<=			16'h80EF;
		end
		32'h00003876: begin
				q			<=			16'h7480;
		end
		32'h00003878: begin
				q			<=			16'h2883;
		end
		32'h0000387A: begin
				q			<=			16'h0401;
		end
		32'h0000387C: begin
				q			<=			16'h1C63;
		end
		32'h0000387E: begin
				q			<=			16'h1805;
		end
		32'h00003880: begin
				q			<=			16'h7A13;
		end
		32'h00003882: begin
				q			<=			16'h001A;
		end
		32'h00003884: begin
				q			<=			16'h0863;
		end
		32'h00003886: begin
				q			<=			16'h180A;
		end
		32'h00003888: begin
				q			<=			16'hC603;
		end
		32'h0000388A: begin
				q			<=			16'h00FA;
		end
		32'h0000388C: begin
				q			<=			16'h2E23;
		end
		32'h0000388E: begin
				q			<=			16'h0BB1;
		end
		32'h00003890: begin
				q			<=			16'h0593;
		end
		32'h00003892: begin
				q			<=			16'h0300;
		end
		32'h00003894: begin
				q			<=			16'h2683;
		end
		32'h00003896: begin
				q			<=			16'h0BC1;
		end
		32'h00003898: begin
				q			<=			16'h8793;
		end
		32'h0000389A: begin
				q			<=			16'hFFF6;
		end
		32'h0000389C: begin
				q			<=			16'h2E23;
		end
		32'h0000389E: begin
				q			<=			16'h0AF1;
		end
		32'h000038A0: begin
				q			<=			16'hC783;
		end
		32'h000038A2: begin
				q			<=			16'hFFF6;
		end
		32'h000038A4: begin
				q			<=			16'h8463;
		end
		32'h000038A6: begin
				q			<=			16'h14C7;
		end
		32'h000038A8: begin
				q			<=			16'h0613;
		end
		32'h000038AA: begin
				q			<=			16'h0390;
		end
		32'h000038AC: begin
				q			<=			16'h9463;
		end
		32'h000038AE: begin
				q			<=			16'h14C7;
		end
		32'h000038B0: begin
				q			<=			16'hC783;
		end
		32'h000038B2: begin
				q			<=			16'h00AA;
		end
		32'h000038B4: begin
				q			<=			16'h8FA3;
		end
		32'h000038B6: begin
				q			<=			16'hFEF6;
		end
		32'h000038B8: begin
				q			<=			16'h8A13;
		end
		32'h000038BA: begin
				q			<=			16'h000D;
		end
		32'h000038BC: begin
				q			<=			16'h0713;
		end
		32'h000038BE: begin
				q			<=			16'h0470;
		end
		32'h000038C0: begin
				q			<=			16'h0A33;
		end
		32'h000038C2: begin
				q			<=			16'h409A;
		end
		32'h000038C4: begin
				q			<=			16'h2C83;
		end
		32'h000038C6: begin
				q			<=			16'h0AC1;
		end
		32'h000038C8: begin
				q			<=			16'h9463;
		end
		32'h000038CA: begin
				q			<=			16'h2AEB;
		end
		32'h000038CC: begin
				q			<=			16'h0713;
		end
		32'h000038CE: begin
				q			<=			16'hFFD0;
		end
		32'h000038D0: begin
				q			<=			16'hC463;
		end
		32'h000038D2: begin
				q			<=			16'h00EC;
		end
		32'h000038D4: begin
				q			<=			16'h5063;
		end
		32'h000038D6: begin
				q			<=			16'h339B;
		end
		32'h000038D8: begin
				q			<=			16'h0D13;
		end
		32'h000038DA: begin
				q			<=			16'hFFED;
		end
		32'h000038DC: begin
				q			<=			16'h8713;
		end
		32'h000038DE: begin
				q			<=			16'hFFFC;
		end
		32'h000038E0: begin
				q			<=			16'h2623;
		end
		32'h000038E2: begin
				q			<=			16'h0AE1;
		end
		32'h000038E4: begin
				q			<=			16'h7613;
		end
		32'h000038E6: begin
				q			<=			16'hFDFD;
		end
		32'h000038E8: begin
				q			<=			16'h0513;
		end
		32'h000038EA: begin
				q			<=			16'h0410;
		end
		32'h000038EC: begin
				q			<=			16'h7693;
		end
		32'h000038EE: begin
				q			<=			16'h0FFD;
		end
		32'h000038F0: begin
				q			<=			16'h0593;
		end
		32'h000038F2: begin
				q			<=			16'h0000;
		end
		32'h000038F4: begin
				q			<=			16'h1863;
		end
		32'h000038F6: begin
				q			<=			16'h00A6;
		end
		32'h000038F8: begin
				q			<=			16'h8693;
		end
		32'h000038FA: begin
				q			<=			16'h00F6;
		end
		32'h000038FC: begin
				q			<=			16'hF693;
		end
		32'h000038FE: begin
				q			<=			16'h0FF6;
		end
		32'h00003900: begin
				q			<=			16'h0593;
		end
		32'h00003902: begin
				q			<=			16'h0010;
		end
		32'h00003904: begin
				q			<=			16'h0A23;
		end
		32'h00003906: begin
				q			<=			16'h0AD1;
		end
		32'h00003908: begin
				q			<=			16'h0793;
		end
		32'h0000390A: begin
				q			<=			16'h02B0;
		end
		32'h0000390C: begin
				q			<=			16'h5863;
		end
		32'h0000390E: begin
				q			<=			16'h0007;
		end
		32'h00003910: begin
				q			<=			16'h0713;
		end
		32'h00003912: begin
				q			<=			16'h0010;
		end
		32'h00003914: begin
				q			<=			16'h0733;
		end
		32'h00003916: begin
				q			<=			16'h4197;
		end
		32'h00003918: begin
				q			<=			16'h0793;
		end
		32'h0000391A: begin
				q			<=			16'h02D0;
		end
		32'h0000391C: begin
				q			<=			16'h0AA3;
		end
		32'h0000391E: begin
				q			<=			16'h0AF1;
		end
		32'h00003920: begin
				q			<=			16'h0793;
		end
		32'h00003922: begin
				q			<=			16'h0090;
		end
		32'h00003924: begin
				q			<=			16'hDA63;
		end
		32'h00003926: begin
				q			<=			16'h28E7;
		end
		32'h00003928: begin
				q			<=			16'h0793;
		end
		32'h0000392A: begin
				q			<=			16'h0C31;
		end
		32'h0000392C: begin
				q			<=			16'h8593;
		end
		32'h0000392E: begin
				q			<=			16'h0007;
		end
		32'h00003930: begin
				q			<=			16'h0513;
		end
		32'h00003932: begin
				q			<=			16'h0090;
		end
		32'h00003934: begin
				q			<=			16'h0813;
		end
		32'h00003936: begin
				q			<=			16'h00A0;
		end
		32'h00003938: begin
				q			<=			16'h66B3;
		end
		32'h0000393A: begin
				q			<=			16'h0307;
		end
		32'h0000393C: begin
				q			<=			16'h8613;
		end
		32'h0000393E: begin
				q			<=			16'hFFF7;
		end
		32'h00003940: begin
				q			<=			16'h4733;
		end
		32'h00003942: begin
				q			<=			16'h0307;
		end
		32'h00003944: begin
				q			<=			16'h8693;
		end
		32'h00003946: begin
				q			<=			16'h0306;
		end
		32'h00003948: begin
				q			<=			16'h8FA3;
		end
		32'h0000394A: begin
				q			<=			16'hFED7;
		end
		32'h0000394C: begin
				q			<=			16'h4863;
		end
		32'h0000394E: begin
				q			<=			16'h24E5;
		end
		32'h00003950: begin
				q			<=			16'h0713;
		end
		32'h00003952: begin
				q			<=			16'h0307;
		end
		32'h00003954: begin
				q			<=			16'h8793;
		end
		32'h00003956: begin
				q			<=			16'hFFE7;
		end
		32'h00003958: begin
				q			<=			16'h0FA3;
		end
		32'h0000395A: begin
				q			<=			16'hFEE6;
		end
		32'h0000395C: begin
				q			<=			16'h0693;
		end
		32'h0000395E: begin
				q			<=			16'h0B61;
		end
		32'h00003960: begin
				q			<=			16'hE263;
		end
		32'h00003962: begin
				q			<=			16'h24B7;
		end
		32'h00003964: begin
				q			<=			16'h0793;
		end
		32'h00003966: begin
				q			<=			16'h0B41;
		end
		32'h00003968: begin
				q			<=			16'h87B3;
		end
		32'h0000396A: begin
				q			<=			16'h40F6;
		end
		32'h0000396C: begin
				q			<=			16'h2823;
		end
		32'h0000396E: begin
				q			<=			16'h02F1;
		end
		32'h00003970: begin
				q			<=			16'h8B33;
		end
		32'h00003972: begin
				q			<=			16'h0147;
		end
		32'h00003974: begin
				q			<=			16'h0793;
		end
		32'h00003976: begin
				q			<=			16'h0010;
		end
		32'h00003978: begin
				q			<=			16'hC663;
		end
		32'h0000397A: begin
				q			<=			16'h0147;
		end
		32'h0000397C: begin
				q			<=			16'h7793;
		end
		32'h0000397E: begin
				q			<=			16'h0014;
		end
		32'h00003980: begin
				q			<=			16'h8663;
		end
		32'h00003982: begin
				q			<=			16'h0007;
		end
		32'h00003984: begin
				q			<=			16'h2783;
		end
		32'h00003986: begin
				q			<=			16'h0141;
		end
		32'h00003988: begin
				q			<=			16'h0B33;
		end
		32'h0000398A: begin
				q			<=			16'h00FB;
		end
		32'h0000398C: begin
				q			<=			16'h7413;
		end
		32'h0000398E: begin
				q			<=			16'hBFF4;
		end
		32'h00003990: begin
				q			<=			16'h6793;
		end
		32'h00003992: begin
				q			<=			16'h1004;
		end
		32'h00003994: begin
				q			<=			16'h2023;
		end
		32'h00003996: begin
				q			<=			16'h02F1;
		end
		32'h00003998: begin
				q			<=			16'h0C13;
		end
		32'h0000399A: begin
				q			<=			16'h0000;
		end
		32'h0000399C: begin
				q			<=			16'h0B93;
		end
		32'h0000399E: begin
				q			<=			16'h0000;
		end
		32'h000039A0: begin
				q			<=			16'h0C93;
		end
		32'h000039A2: begin
				q			<=			16'h0000;
		end
		32'h000039A4: begin
				q			<=			16'h2783;
		end
		32'h000039A6: begin
				q			<=			16'h0381;
		end
		32'h000039A8: begin
				q			<=			16'h8663;
		end
		32'h000039AA: begin
				q			<=			16'h0007;
		end
		32'h000039AC: begin
				q			<=			16'h0713;
		end
		32'h000039AE: begin
				q			<=			16'h02D0;
		end
		32'h000039B0: begin
				q			<=			16'h03A3;
		end
		32'h000039B2: begin
				q			<=			16'h0AE1;
		end
		32'h000039B4: begin
				q			<=			16'h2403;
		end
		32'h000039B6: begin
				q			<=			16'h0201;
		end
		32'h000039B8: begin
				q			<=			16'h0D93;
		end
		32'h000039BA: begin
				q			<=			16'h0000;
		end
		32'h000039BC: begin
				q			<=			16'h006F;
		end
		32'h000039BE: begin
				q			<=			16'h4880;
		end
		32'h000039C0: begin
				q			<=			16'h2223;
		end
		32'h000039C2: begin
				q			<=			16'h0001;
		end
		32'h000039C4: begin
				q			<=			16'h0493;
		end
		32'h000039C6: begin
				q			<=			16'h12C1;
		end
		32'h000039C8: begin
				q			<=			16'hF06F;
		end
		32'h000039CA: begin
				q			<=			16'hB9DF;
		end
		32'h000039CC: begin
				q			<=			16'h2223;
		end
		32'h000039CE: begin
				q			<=			16'h00A1;
		end
		32'h000039D0: begin
				q			<=			16'hF06F;
		end
		32'h000039D2: begin
				q			<=			16'hB95F;
		end
		32'h000039D4: begin
				q			<=			16'h2223;
		end
		32'h000039D6: begin
				q			<=			16'h0001;
		end
		32'h000039D8: begin
				q			<=			16'h0B13;
		end
		32'h000039DA: begin
				q			<=			16'h0060;
		end
		32'h000039DC: begin
				q			<=			16'hF06F;
		end
		32'h000039DE: begin
				q			<=			16'hB89F;
		end
		32'h000039E0: begin
				q			<=			16'h2223;
		end
		32'h000039E2: begin
				q			<=			16'h0161;
		end
		32'h000039E4: begin
				q			<=			16'h0B13;
		end
		32'h000039E6: begin
				q			<=			16'h0010;
		end
		32'h000039E8: begin
				q			<=			16'hF06F;
		end
		32'h000039EA: begin
				q			<=			16'hB7DF;
		end
		32'h000039EC: begin
				q			<=			16'h8FA3;
		end
		32'h000039EE: begin
				q			<=			16'hFEB6;
		end
		32'h000039F0: begin
				q			<=			16'hF06F;
		end
		32'h000039F2: begin
				q			<=			16'hEA5F;
		end
		32'h000039F4: begin
				q			<=			16'h8793;
		end
		32'h000039F6: begin
				q			<=			16'h0017;
		end
		32'h000039F8: begin
				q			<=			16'hF793;
		end
		32'h000039FA: begin
				q			<=			16'h0FF7;
		end
		32'h000039FC: begin
				q			<=			16'hF06F;
		end
		32'h000039FE: begin
				q			<=			16'hEB9F;
		end
		32'h00003A00: begin
				q			<=			16'h0A13;
		end
		32'h00003A02: begin
				q			<=			16'h001A;
		end
		32'h00003A04: begin
				q			<=			16'h0FA3;
		end
		32'h00003A06: begin
				q			<=			16'hFEEA;
		end
		32'h00003A08: begin
				q			<=			16'h07B3;
		end
		32'h00003A0A: begin
				q			<=			16'h414C;
		end
		32'h00003A0C: begin
				q			<=			16'hDAE3;
		end
		32'h00003A0E: begin
				q			<=			16'hFE07;
		end
		32'h00003A10: begin
				q			<=			16'hF06F;
		end
		32'h00003A12: begin
				q			<=			16'hEADF;
		end
		32'h00003A14: begin
				q			<=			16'h2783;
		end
		32'h00003A16: begin
				q			<=			16'h03C1;
		end
		32'h00003A18: begin
				q			<=			16'h8A13;
		end
		32'h00003A1A: begin
				q			<=			16'h000D;
		end
		32'h00003A1C: begin
				q			<=			16'h0713;
		end
		32'h00003A1E: begin
				q			<=			16'h0300;
		end
		32'h00003A20: begin
				q			<=			16'h8C33;
		end
		32'h00003A22: begin
				q			<=			16'h00FD;
		end
		32'h00003A24: begin
				q			<=			16'hF06F;
		end
		32'h00003A26: begin
				q			<=			16'hFE5F;
		end
		32'h00003A28: begin
				q			<=			16'h0793;
		end
		32'h00003A2A: begin
				q			<=			16'h0460;
		end
		32'h00003A2C: begin
				q			<=			16'h8E63;
		end
		32'h00003A2E: begin
				q			<=			16'h00FB;
		end
		32'h00003A30: begin
				q			<=			16'h0793;
		end
		32'h00003A32: begin
				q			<=			16'h0450;
		end
		32'h00003A34: begin
				q			<=			16'h0C13;
		end
		32'h00003A36: begin
				q			<=			16'h001B;
		end
		32'h00003A38: begin
				q			<=			16'h8463;
		end
		32'h00003A3A: begin
				q			<=			16'h00FB;
		end
		32'h00003A3C: begin
				q			<=			16'h0C13;
		end
		32'h00003A3E: begin
				q			<=			16'h000B;
		end
		32'h00003A40: begin
				q			<=			16'h0613;
		end
		32'h00003A42: begin
				q			<=			16'h0020;
		end
		32'h00003A44: begin
				q			<=			16'h006F;
		end
		32'h00003A46: begin
				q			<=			16'h00C0;
		end
		32'h00003A48: begin
				q			<=			16'h0C13;
		end
		32'h00003A4A: begin
				q			<=			16'h000B;
		end
		32'h00003A4C: begin
				q			<=			16'h0613;
		end
		32'h00003A4E: begin
				q			<=			16'h0030;
		end
		32'h00003A50: begin
				q			<=			16'h0793;
		end
		32'h00003A52: begin
				q			<=			16'h0B01;
		end
		32'h00003A54: begin
				q			<=			16'h0813;
		end
		32'h00003A56: begin
				q			<=			16'h0BC1;
		end
		32'h00003A58: begin
				q			<=			16'h0713;
		end
		32'h00003A5A: begin
				q			<=			16'h0AC1;
		end
		32'h00003A5C: begin
				q			<=			16'h0693;
		end
		32'h00003A5E: begin
				q			<=			16'h000C;
		end
		32'h00003A60: begin
				q			<=			16'h0593;
		end
		32'h00003A62: begin
				q			<=			16'h0901;
		end
		32'h00003A64: begin
				q			<=			16'h0513;
		end
		32'h00003A66: begin
				q			<=			16'h0009;
		end
		32'h00003A68: begin
				q			<=			16'h2023;
		end
		32'h00003A6A: begin
				q			<=			16'h0511;
		end
		32'h00003A6C: begin
				q			<=			16'h2823;
		end
		32'h00003A6E: begin
				q			<=			16'h09C1;
		end
		32'h00003A70: begin
				q			<=			16'h2E23;
		end
		32'h00003A72: begin
				q			<=			16'h03C1;
		end
		32'h00003A74: begin
				q			<=			16'h2A23;
		end
		32'h00003A76: begin
				q			<=			16'h09B1;
		end
		32'h00003A78: begin
				q			<=			16'h2C23;
		end
		32'h00003A7A: begin
				q			<=			16'h0991;
		end
		32'h00003A7C: begin
				q			<=			16'h2E23;
		end
		32'h00003A7E: begin
				q			<=			16'h0951;
		end
		32'h00003A80: begin
				q			<=			16'h3097;
		end
		32'h00003A82: begin
				q			<=			16'h0000;
		end
		32'h00003A84: begin
				q			<=			16'h80E7;
		end
		32'h00003A86: begin
				q			<=			16'hB980;
		end
		32'h00003A88: begin
				q			<=			16'h0793;
		end
		32'h00003A8A: begin
				q			<=			16'h0470;
		end
		32'h00003A8C: begin
				q			<=			16'h0493;
		end
		32'h00003A8E: begin
				q			<=			16'h0005;
		end
		32'h00003A90: begin
				q			<=			16'h2E03;
		end
		32'h00003A92: begin
				q			<=			16'h03C1;
		end
		32'h00003A94: begin
				q			<=			16'h2883;
		end
		32'h00003A96: begin
				q			<=			16'h0401;
		end
		32'h00003A98: begin
				q			<=			16'h9663;
		end
		32'h00003A9A: begin
				q			<=			16'h00FB;
		end
		32'h00003A9C: begin
				q			<=			16'h7793;
		end
		32'h00003A9E: begin
				q			<=			16'h0014;
		end
		32'h00003AA0: begin
				q			<=			16'h8863;
		end
		32'h00003AA2: begin
				q			<=			16'h0A07;
		end
		32'h00003AA4: begin
				q			<=			16'h0793;
		end
		32'h00003AA6: begin
				q			<=			16'h0460;
		end
		32'h00003AA8: begin
				q			<=			16'h8A33;
		end
		32'h00003AAA: begin
				q			<=			16'h0184;
		end
		32'h00003AAC: begin
				q			<=			16'h9263;
		end
		32'h00003AAE: begin
				q			<=			16'h06FB;
		end
		32'h00003AB0: begin
				q			<=			16'hC703;
		end
		32'h00003AB2: begin
				q			<=			16'h0004;
		end
		32'h00003AB4: begin
				q			<=			16'h0793;
		end
		32'h00003AB6: begin
				q			<=			16'h0300;
		end
		32'h00003AB8: begin
				q			<=			16'h1863;
		end
		32'h00003ABA: begin
				q			<=			16'h04F7;
		end
		32'h00003ABC: begin
				q			<=			16'h0593;
		end
		32'h00003ABE: begin
				q			<=			16'h0801;
		end
		32'h00003AC0: begin
				q			<=			16'h0513;
		end
		32'h00003AC2: begin
				q			<=			16'h0901;
		end
		32'h00003AC4: begin
				q			<=			16'h2023;
		end
		32'h00003AC6: begin
				q			<=			16'h0511;
		end
		32'h00003AC8: begin
				q			<=			16'h2823;
		end
		32'h00003ACA: begin
				q			<=			16'h09C1;
		end
		32'h00003ACC: begin
				q			<=			16'h2E23;
		end
		32'h00003ACE: begin
				q			<=			16'h03C1;
		end
		32'h00003AD0: begin
				q			<=			16'h2A23;
		end
		32'h00003AD2: begin
				q			<=			16'h09B1;
		end
		32'h00003AD4: begin
				q			<=			16'h2C23;
		end
		32'h00003AD6: begin
				q			<=			16'h0991;
		end
		32'h00003AD8: begin
				q			<=			16'h2E23;
		end
		32'h00003ADA: begin
				q			<=			16'h0951;
		end
		32'h00003ADC: begin
				q			<=			16'h2023;
		end
		32'h00003ADE: begin
				q			<=			16'h0801;
		end
		32'h00003AE0: begin
				q			<=			16'h2223;
		end
		32'h00003AE2: begin
				q			<=			16'h0801;
		end
		32'h00003AE4: begin
				q			<=			16'h2423;
		end
		32'h00003AE6: begin
				q			<=			16'h0801;
		end
		32'h00003AE8: begin
				q			<=			16'h2623;
		end
		32'h00003AEA: begin
				q			<=			16'h0801;
		end
		32'h00003AEC: begin
				q			<=			16'h80EF;
		end
		32'h00003AEE: begin
				q			<=			16'h4D00;
		end
		32'h00003AF0: begin
				q			<=			16'h2E03;
		end
		32'h00003AF2: begin
				q			<=			16'h03C1;
		end
		32'h00003AF4: begin
				q			<=			16'h2883;
		end
		32'h00003AF6: begin
				q			<=			16'h0401;
		end
		32'h00003AF8: begin
				q			<=			16'h0863;
		end
		32'h00003AFA: begin
				q			<=			16'h0005;
		end
		32'h00003AFC: begin
				q			<=			16'h0793;
		end
		32'h00003AFE: begin
				q			<=			16'h0010;
		end
		32'h00003B00: begin
				q			<=			16'h8C33;
		end
		32'h00003B02: begin
				q			<=			16'h4187;
		end
		32'h00003B04: begin
				q			<=			16'h2623;
		end
		32'h00003B06: begin
				q			<=			16'h0B81;
		end
		32'h00003B08: begin
				q			<=			16'h2783;
		end
		32'h00003B0A: begin
				q			<=			16'h0AC1;
		end
		32'h00003B0C: begin
				q			<=			16'h0A33;
		end
		32'h00003B0E: begin
				q			<=			16'h00FA;
		end
		32'h00003B10: begin
				q			<=			16'h0593;
		end
		32'h00003B12: begin
				q			<=			16'h0801;
		end
		32'h00003B14: begin
				q			<=			16'h0513;
		end
		32'h00003B16: begin
				q			<=			16'h0901;
		end
		32'h00003B18: begin
				q			<=			16'h2E23;
		end
		32'h00003B1A: begin
				q			<=			16'h0311;
		end
		32'h00003B1C: begin
				q			<=			16'h2823;
		end
		32'h00003B1E: begin
				q			<=			16'h09C1;
		end
		32'h00003B20: begin
				q			<=			16'h2A23;
		end
		32'h00003B22: begin
				q			<=			16'h09B1;
		end
		32'h00003B24: begin
				q			<=			16'h2C23;
		end
		32'h00003B26: begin
				q			<=			16'h0991;
		end
		32'h00003B28: begin
				q			<=			16'h2E23;
		end
		32'h00003B2A: begin
				q			<=			16'h0951;
		end
		32'h00003B2C: begin
				q			<=			16'h2023;
		end
		32'h00003B2E: begin
				q			<=			16'h0801;
		end
		32'h00003B30: begin
				q			<=			16'h2223;
		end
		32'h00003B32: begin
				q			<=			16'h0801;
		end
		32'h00003B34: begin
				q			<=			16'h2423;
		end
		32'h00003B36: begin
				q			<=			16'h0801;
		end
		32'h00003B38: begin
				q			<=			16'h2623;
		end
		32'h00003B3A: begin
				q			<=			16'h0801;
		end
		32'h00003B3C: begin
				q			<=			16'h80EF;
		end
		32'h00003B3E: begin
				q			<=			16'h4800;
		end
		32'h00003B40: begin
				q			<=			16'h2883;
		end
		32'h00003B42: begin
				q			<=			16'h03C1;
		end
		32'h00003B44: begin
				q			<=			16'h0713;
		end
		32'h00003B46: begin
				q			<=			16'h0300;
		end
		32'h00003B48: begin
				q			<=			16'h1E63;
		end
		32'h00003B4A: begin
				q			<=			16'h0005;
		end
		32'h00003B4C: begin
				q			<=			16'h2E23;
		end
		32'h00003B4E: begin
				q			<=			16'h0B41;
		end
		32'h00003B50: begin
				q			<=			16'h2A03;
		end
		32'h00003B52: begin
				q			<=			16'h0BC1;
		end
		32'h00003B54: begin
				q			<=			16'hF06F;
		end
		32'h00003B56: begin
				q			<=			16'hD69F;
		end
		32'h00003B58: begin
				q			<=			16'h8693;
		end
		32'h00003B5A: begin
				q			<=			16'h0017;
		end
		32'h00003B5C: begin
				q			<=			16'h2E23;
		end
		32'h00003B5E: begin
				q			<=			16'h0AD1;
		end
		32'h00003B60: begin
				q			<=			16'h8023;
		end
		32'h00003B62: begin
				q			<=			16'h00E7;
		end
		32'h00003B64: begin
				q			<=			16'h2783;
		end
		32'h00003B66: begin
				q			<=			16'h0BC1;
		end
		32'h00003B68: begin
				q			<=			16'hE8E3;
		end
		32'h00003B6A: begin
				q			<=			16'hFF47;
		end
		32'h00003B6C: begin
				q			<=			16'hF06F;
		end
		32'h00003B6E: begin
				q			<=			16'hFE5F;
		end
		32'h00003B70: begin
				q			<=			16'h0713;
		end
		32'h00003B72: begin
				q			<=			16'h0460;
		end
		32'h00003B74: begin
				q			<=			16'h94E3;
		end
		32'h00003B76: begin
				q			<=			16'hD6EB;
		end
		32'h00003B78: begin
				q			<=			16'h5263;
		end
		32'h00003B7A: begin
				q			<=			16'h0790;
		end
		32'h00003B7C: begin
				q			<=			16'h1663;
		end
		32'h00003B7E: begin
				q			<=			16'h000B;
		end
		32'h00003B80: begin
				q			<=			16'h7713;
		end
		32'h00003B82: begin
				q			<=			16'h0014;
		end
		32'h00003B84: begin
				q			<=			16'h0263;
		end
		32'h00003B86: begin
				q			<=			16'h0C07;
		end
		32'h00003B88: begin
				q			<=			16'h2783;
		end
		32'h00003B8A: begin
				q			<=			16'h0141;
		end
		32'h00003B8C: begin
				q			<=			16'h8733;
		end
		32'h00003B8E: begin
				q			<=			16'h00FC;
		end
		32'h00003B90: begin
				q			<=			16'h0B33;
		end
		32'h00003B92: begin
				q			<=			16'h00EB;
		end
		32'h00003B94: begin
				q			<=			16'h0D13;
		end
		32'h00003B96: begin
				q			<=			16'h0660;
		end
		32'h00003B98: begin
				q			<=			16'h006F;
		end
		32'h00003B9A: begin
				q			<=			16'h0940;
		end
		32'h00003B9C: begin
				q			<=			16'h0793;
		end
		32'h00003B9E: begin
				q			<=			16'h0006;
		end
		32'h00003BA0: begin
				q			<=			16'hF06F;
		end
		32'h00003BA2: begin
				q			<=			16'hD95F;
		end
		32'h00003BA4: begin
				q			<=			16'h8793;
		end
		32'h00003BA6: begin
				q			<=			16'h0017;
		end
		32'h00003BA8: begin
				q			<=			16'hC703;
		end
		32'h00003BAA: begin
				q			<=			16'hFFF7;
		end
		32'h00003BAC: begin
				q			<=			16'h8693;
		end
		32'h00003BAE: begin
				q			<=			16'h0016;
		end
		32'h00003BB0: begin
				q			<=			16'h8FA3;
		end
		32'h00003BB2: begin
				q			<=			16'hFEE6;
		end
		32'h00003BB4: begin
				q			<=			16'hF06F;
		end
		32'h00003BB6: begin
				q			<=			16'hDADF;
		end
		32'h00003BB8: begin
				q			<=			16'h0793;
		end
		32'h00003BBA: begin
				q			<=			16'h0B61;
		end
		32'h00003BBC: begin
				q			<=			16'h9863;
		end
		32'h00003BBE: begin
				q			<=			16'h0005;
		end
		32'h00003BC0: begin
				q			<=			16'h0793;
		end
		32'h00003BC2: begin
				q			<=			16'h0300;
		end
		32'h00003BC4: begin
				q			<=			16'h0B23;
		end
		32'h00003BC6: begin
				q			<=			16'h0AF1;
		end
		32'h00003BC8: begin
				q			<=			16'h0793;
		end
		32'h00003BCA: begin
				q			<=			16'h0B71;
		end
		32'h00003BCC: begin
				q			<=			16'h0713;
		end
		32'h00003BCE: begin
				q			<=			16'h0307;
		end
		32'h00003BD0: begin
				q			<=			16'h8693;
		end
		32'h00003BD2: begin
				q			<=			16'h0017;
		end
		32'h00003BD4: begin
				q			<=			16'h8023;
		end
		32'h00003BD6: begin
				q			<=			16'h00E7;
		end
		32'h00003BD8: begin
				q			<=			16'hF06F;
		end
		32'h00003BDA: begin
				q			<=			16'hD8DF;
		end
		32'h00003BDC: begin
				q			<=			16'h1663;
		end
		32'h00003BDE: begin
				q			<=			16'h000B;
		end
		32'h00003BE0: begin
				q			<=			16'h7713;
		end
		32'h00003BE2: begin
				q			<=			16'h0014;
		end
		32'h00003BE4: begin
				q			<=			16'h0663;
		end
		32'h00003BE6: begin
				q			<=			16'h0607;
		end
		32'h00003BE8: begin
				q			<=			16'h2783;
		end
		32'h00003BEA: begin
				q			<=			16'h0141;
		end
		32'h00003BEC: begin
				q			<=			16'h8713;
		end
		32'h00003BEE: begin
				q			<=			16'h0017;
		end
		32'h00003BF0: begin
				q			<=			16'hF06F;
		end
		32'h00003BF2: begin
				q			<=			16'hFA1F;
		end
		32'h00003BF4: begin
				q			<=			16'hC063;
		end
		32'h00003BF6: begin
				q			<=			16'h034C;
		end
		32'h00003BF8: begin
				q			<=			16'h7713;
		end
		32'h00003BFA: begin
				q			<=			16'h0014;
		end
		32'h00003BFC: begin
				q			<=			16'h8B13;
		end
		32'h00003BFE: begin
				q			<=			16'h000C;
		end
		32'h00003C00: begin
				q			<=			16'h0663;
		end
		32'h00003C02: begin
				q			<=			16'h0007;
		end
		32'h00003C04: begin
				q			<=			16'h2783;
		end
		32'h00003C06: begin
				q			<=			16'h0141;
		end
		32'h00003C08: begin
				q			<=			16'h8B33;
		end
		32'h00003C0A: begin
				q			<=			16'h00FC;
		end
		32'h00003C0C: begin
				q			<=			16'h0D13;
		end
		32'h00003C0E: begin
				q			<=			16'h0670;
		end
		32'h00003C10: begin
				q			<=			16'h006F;
		end
		32'h00003C12: begin
				q			<=			16'h01C0;
		end
		32'h00003C14: begin
				q			<=			16'h2783;
		end
		32'h00003C16: begin
				q			<=			16'h0141;
		end
		32'h00003C18: begin
				q			<=			16'h0D13;
		end
		32'h00003C1A: begin
				q			<=			16'h0670;
		end
		32'h00003C1C: begin
				q			<=			16'h0B33;
		end
		32'h00003C1E: begin
				q			<=			16'h00FA;
		end
		32'h00003C20: begin
				q			<=			16'h4663;
		end
		32'h00003C22: begin
				q			<=			16'h0190;
		end
		32'h00003C24: begin
				q			<=			16'h0333;
		end
		32'h00003C26: begin
				q			<=			16'h419B;
		end
		32'h00003C28: begin
				q			<=			16'h0B13;
		end
		32'h00003C2A: begin
				q			<=			16'h0013;
		end
		32'h00003C2C: begin
				q			<=			16'h7B93;
		end
		32'h00003C2E: begin
				q			<=			16'h4004;
		end
		32'h00003C30: begin
				q			<=			16'h0C13;
		end
		32'h00003C32: begin
				q			<=			16'h0000;
		end
		32'h00003C34: begin
				q			<=			16'h88E3;
		end
		32'h00003C36: begin
				q			<=			16'hD60B;
		end
		32'h00003C38: begin
				q			<=			16'h0B93;
		end
		32'h00003C3A: begin
				q			<=			16'h0000;
		end
		32'h00003C3C: begin
				q			<=			16'h54E3;
		end
		32'h00003C3E: begin
				q			<=			16'hD790;
		end
		32'h00003C40: begin
				q			<=			16'h0693;
		end
		32'h00003C42: begin
				q			<=			16'h0FF0;
		end
		32'h00003C44: begin
				q			<=			16'h006F;
		end
		32'h00003C46: begin
				q			<=			16'h0380;
		end
		32'h00003C48: begin
				q			<=			16'h8B13;
		end
		32'h00003C4A: begin
				q			<=			16'h000C;
		end
		32'h00003C4C: begin
				q			<=			16'hF06F;
		end
		32'h00003C4E: begin
				q			<=			16'hF49F;
		end
		32'h00003C50: begin
				q			<=			16'h0D13;
		end
		32'h00003C52: begin
				q			<=			16'h0660;
		end
		32'h00003C54: begin
				q			<=			16'h0B13;
		end
		32'h00003C56: begin
				q			<=			16'h0010;
		end
		32'h00003C58: begin
				q			<=			16'hF06F;
		end
		32'h00003C5A: begin
				q			<=			16'hFD5F;
		end
		32'h00003C5C: begin
				q			<=			16'h5663;
		end
		32'h00003C5E: begin
				q			<=			16'h0397;
		end
		32'h00003C60: begin
				q			<=			16'h2783;
		end
		32'h00003C62: begin
				q			<=			16'h0081;
		end
		32'h00003C64: begin
				q			<=			16'h8CB3;
		end
		32'h00003C66: begin
				q			<=			16'h40EC;
		end
		32'h00003C68: begin
				q			<=			16'hC703;
		end
		32'h00003C6A: begin
				q			<=			16'h0017;
		end
		32'h00003C6C: begin
				q			<=			16'h0863;
		end
		32'h00003C6E: begin
				q			<=			16'h0207;
		end
		32'h00003C70: begin
				q			<=			16'h8793;
		end
		32'h00003C72: begin
				q			<=			16'h0017;
		end
		32'h00003C74: begin
				q			<=			16'h8B93;
		end
		32'h00003C76: begin
				q			<=			16'h001B;
		end
		32'h00003C78: begin
				q			<=			16'h2423;
		end
		32'h00003C7A: begin
				q			<=			16'h00F1;
		end
		32'h00003C7C: begin
				q			<=			16'h2783;
		end
		32'h00003C7E: begin
				q			<=			16'h0081;
		end
		32'h00003C80: begin
				q			<=			16'hC703;
		end
		32'h00003C82: begin
				q			<=			16'h0007;
		end
		32'h00003C84: begin
				q			<=			16'h1CE3;
		end
		32'h00003C86: begin
				q			<=			16'hFCD7;
		end
		32'h00003C88: begin
				q			<=			16'h2783;
		end
		32'h00003C8A: begin
				q			<=			16'h0241;
		end
		32'h00003C8C: begin
				q			<=			16'h8733;
		end
		32'h00003C8E: begin
				q			<=			16'h018B;
		end
		32'h00003C90: begin
				q			<=			16'h0733;
		end
		32'h00003C92: begin
				q			<=			16'h02F7;
		end
		32'h00003C94: begin
				q			<=			16'h0B33;
		end
		32'h00003C96: begin
				q			<=			16'h0167;
		end
		32'h00003C98: begin
				q			<=			16'hF06F;
		end
		32'h00003C9A: begin
				q			<=			16'hD0DF;
		end
		32'h00003C9C: begin
				q			<=			16'h0C13;
		end
		32'h00003C9E: begin
				q			<=			16'h001C;
		end
		32'h00003CA0: begin
				q			<=			16'hF06F;
		end
		32'h00003CA2: begin
				q			<=			16'hFDDF;
		end
		32'h00003CA4: begin
				q			<=			16'h8713;
		end
		32'h00003CA6: begin
				q			<=			16'h004A;
		end
		32'h00003CA8: begin
				q			<=			16'h2623;
		end
		32'h00003CAA: begin
				q			<=			16'h00E1;
		end
		32'h00003CAC: begin
				q			<=			16'h7713;
		end
		32'h00003CAE: begin
				q			<=			16'h0204;
		end
		32'h00003CB0: begin
				q			<=			16'hA783;
		end
		32'h00003CB2: begin
				q			<=			16'h000A;
		end
		32'h00003CB4: begin
				q			<=			16'h0063;
		end
		32'h00003CB6: begin
				q			<=			16'h0207;
		end
		32'h00003CB8: begin
				q			<=			16'h2703;
		end
		32'h00003CBA: begin
				q			<=			16'h0181;
		end
		32'h00003CBC: begin
				q			<=			16'hA023;
		end
		32'h00003CBE: begin
				q			<=			16'h00E7;
		end
		32'h00003CC0: begin
				q			<=			16'h5713;
		end
		32'h00003CC2: begin
				q			<=			16'h41F7;
		end
		32'h00003CC4: begin
				q			<=			16'hA223;
		end
		32'h00003CC6: begin
				q			<=			16'h00E7;
		end
		32'h00003CC8: begin
				q			<=			16'h2A83;
		end
		32'h00003CCA: begin
				q			<=			16'h00C1;
		end
		32'h00003CCC: begin
				q			<=			16'h2483;
		end
		32'h00003CCE: begin
				q			<=			16'h0101;
		end
		32'h00003CD0: begin
				q			<=			16'hF06F;
		end
		32'h00003CD2: begin
				q			<=			16'hAF0F;
		end
		32'h00003CD4: begin
				q			<=			16'h7713;
		end
		32'h00003CD6: begin
				q			<=			16'h0104;
		end
		32'h00003CD8: begin
				q			<=			16'h0863;
		end
		32'h00003CDA: begin
				q			<=			16'h0007;
		end
		32'h00003CDC: begin
				q			<=			16'h2703;
		end
		32'h00003CDE: begin
				q			<=			16'h0181;
		end
		32'h00003CE0: begin
				q			<=			16'hA023;
		end
		32'h00003CE2: begin
				q			<=			16'h00E7;
		end
		32'h00003CE4: begin
				q			<=			16'hF06F;
		end
		32'h00003CE6: begin
				q			<=			16'hFE5F;
		end
		32'h00003CE8: begin
				q			<=			16'h7713;
		end
		32'h00003CEA: begin
				q			<=			16'h0404;
		end
		32'h00003CEC: begin
				q			<=			16'h0863;
		end
		32'h00003CEE: begin
				q			<=			16'h0007;
		end
		32'h00003CF0: begin
				q			<=			16'h5703;
		end
		32'h00003CF2: begin
				q			<=			16'h0181;
		end
		32'h00003CF4: begin
				q			<=			16'h9023;
		end
		32'h00003CF6: begin
				q			<=			16'h00E7;
		end
		32'h00003CF8: begin
				q			<=			16'hF06F;
		end
		32'h00003CFA: begin
				q			<=			16'hFD1F;
		end
		32'h00003CFC: begin
				q			<=			16'h7413;
		end
		32'h00003CFE: begin
				q			<=			16'h2004;
		end
		32'h00003D00: begin
				q			<=			16'h0EE3;
		end
		32'h00003D02: begin
				q			<=			16'hFC04;
		end
		32'h00003D04: begin
				q			<=			16'h4703;
		end
		32'h00003D06: begin
				q			<=			16'h0181;
		end
		32'h00003D08: begin
				q			<=			16'h8023;
		end
		32'h00003D0A: begin
				q			<=			16'h00E7;
		end
		32'h00003D0C: begin
				q			<=			16'hF06F;
		end
		32'h00003D0E: begin
				q			<=			16'hFBDF;
		end
		32'h00003D10: begin
				q			<=			16'h6413;
		end
		32'h00003D12: begin
				q			<=			16'h0104;
		end
		32'h00003D14: begin
				q			<=			16'h7793;
		end
		32'h00003D16: begin
				q			<=			16'h0204;
		end
		32'h00003D18: begin
				q			<=			16'h8863;
		end
		32'h00003D1A: begin
				q			<=			16'h0407;
		end
		32'h00003D1C: begin
				q			<=			16'h8A93;
		end
		32'h00003D1E: begin
				q			<=			16'h007A;
		end
		32'h00003D20: begin
				q			<=			16'hFA93;
		end
		32'h00003D22: begin
				q			<=			16'hFF8A;
		end
		32'h00003D24: begin
				q			<=			16'hAC03;
		end
		32'h00003D26: begin
				q			<=			16'h000A;
		end
		32'h00003D28: begin
				q			<=			16'hAC83;
		end
		32'h00003D2A: begin
				q			<=			16'h004A;
		end
		32'h00003D2C: begin
				q			<=			16'h8793;
		end
		32'h00003D2E: begin
				q			<=			16'h008A;
		end
		32'h00003D30: begin
				q			<=			16'h2623;
		end
		32'h00003D32: begin
				q			<=			16'h00F1;
		end
		32'h00003D34: begin
				q			<=			16'h7413;
		end
		32'h00003D36: begin
				q			<=			16'hBFF4;
		end
		32'h00003D38: begin
				q			<=			16'h0793;
		end
		32'h00003D3A: begin
				q			<=			16'h0000;
		end
		32'h00003D3C: begin
				q			<=			16'h03A3;
		end
		32'h00003D3E: begin
				q			<=			16'h0A01;
		end
		32'h00003D40: begin
				q			<=			16'h0713;
		end
		32'h00003D42: begin
				q			<=			16'hFFF0;
		end
		32'h00003D44: begin
				q			<=			16'h0C63;
		end
		32'h00003D46: begin
				q			<=			16'h42EB;
		end
		32'h00003D48: begin
				q			<=			16'h0713;
		end
		32'h00003D4A: begin
				q			<=			16'h0004;
		end
		32'h00003D4C: begin
				q			<=			16'h66B3;
		end
		32'h00003D4E: begin
				q			<=			16'h019C;
		end
		32'h00003D50: begin
				q			<=			16'h7413;
		end
		32'h00003D52: begin
				q			<=			16'hF7F4;
		end
		32'h00003D54: begin
				q			<=			16'h9463;
		end
		32'h00003D56: begin
				q			<=			16'h4206;
		end
		32'h00003D58: begin
				q			<=			16'h0263;
		end
		32'h00003D5A: begin
				q			<=			16'h5A0B;
		end
		32'h00003D5C: begin
				q			<=			16'h0713;
		end
		32'h00003D5E: begin
				q			<=			16'h0010;
		end
		32'h00003D60: begin
				q			<=			16'h9263;
		end
		32'h00003D62: begin
				q			<=			16'h42E7;
		end
		32'h00003D64: begin
				q			<=			16'hF06F;
		end
		32'h00003D66: begin
				q			<=			16'hDB0F;
		end
		32'h00003D68: begin
				q			<=			16'h8793;
		end
		32'h00003D6A: begin
				q			<=			16'h004A;
		end
		32'h00003D6C: begin
				q			<=			16'h2623;
		end
		32'h00003D6E: begin
				q			<=			16'h00F1;
		end
		32'h00003D70: begin
				q			<=			16'h7793;
		end
		32'h00003D72: begin
				q			<=			16'h0104;
		end
		32'h00003D74: begin
				q			<=			16'h8663;
		end
		32'h00003D76: begin
				q			<=			16'h0007;
		end
		32'h00003D78: begin
				q			<=			16'hAC03;
		end
		32'h00003D7A: begin
				q			<=			16'h000A;
		end
		32'h00003D7C: begin
				q			<=			16'h006F;
		end
		32'h00003D7E: begin
				q			<=			16'h0100;
		end
		32'h00003D80: begin
				q			<=			16'h7793;
		end
		32'h00003D82: begin
				q			<=			16'h0404;
		end
		32'h00003D84: begin
				q			<=			16'h8863;
		end
		32'h00003D86: begin
				q			<=			16'h0007;
		end
		32'h00003D88: begin
				q			<=			16'hDC03;
		end
		32'h00003D8A: begin
				q			<=			16'h000A;
		end
		32'h00003D8C: begin
				q			<=			16'h0C93;
		end
		32'h00003D8E: begin
				q			<=			16'h0000;
		end
		32'h00003D90: begin
				q			<=			16'hF06F;
		end
		32'h00003D92: begin
				q			<=			16'hFA5F;
		end
		32'h00003D94: begin
				q			<=			16'h7793;
		end
		32'h00003D96: begin
				q			<=			16'h2004;
		end
		32'h00003D98: begin
				q			<=			16'h80E3;
		end
		32'h00003D9A: begin
				q			<=			16'hFE07;
		end
		32'h00003D9C: begin
				q			<=			16'hCC03;
		end
		32'h00003D9E: begin
				q			<=			16'h000A;
		end
		32'h00003DA0: begin
				q			<=			16'hF06F;
		end
		32'h00003DA2: begin
				q			<=			16'hFEDF;
		end
		32'h00003DA4: begin
				q			<=			16'h8793;
		end
		32'h00003DA6: begin
				q			<=			16'h004A;
		end
		32'h00003DA8: begin
				q			<=			16'h2623;
		end
		32'h00003DAA: begin
				q			<=			16'h00F1;
		end
		32'h00003DAC: begin
				q			<=			16'h87B7;
		end
		32'h00003DAE: begin
				q			<=			16'hFFFF;
		end
		32'h00003DB0: begin
				q			<=			16'hC793;
		end
		32'h00003DB2: begin
				q			<=			16'h8307;
		end
		32'h00003DB4: begin
				q			<=			16'h1423;
		end
		32'h00003DB6: begin
				q			<=			16'h0AF1;
		end
		32'h00003DB8: begin
				q			<=			16'hC797;
		end
		32'h00003DBA: begin
				q			<=			16'h0000;
		end
		32'h00003DBC: begin
				q			<=			16'h8793;
		end
		32'h00003DBE: begin
				q			<=			16'hFCC7;
		end
		32'h00003DC0: begin
				q			<=			16'h2A23;
		end
		32'h00003DC2: begin
				q			<=			16'h02F1;
		end
		32'h00003DC4: begin
				q			<=			16'hAC03;
		end
		32'h00003DC6: begin
				q			<=			16'h000A;
		end
		32'h00003DC8: begin
				q			<=			16'h0C93;
		end
		32'h00003DCA: begin
				q			<=			16'h0000;
		end
		32'h00003DCC: begin
				q			<=			16'h6413;
		end
		32'h00003DCE: begin
				q			<=			16'h0024;
		end
		32'h00003DD0: begin
				q			<=			16'h0793;
		end
		32'h00003DD2: begin
				q			<=			16'h0020;
		end
		32'h00003DD4: begin
				q			<=			16'h0D13;
		end
		32'h00003DD6: begin
				q			<=			16'h0780;
		end
		32'h00003DD8: begin
				q			<=			16'hF06F;
		end
		32'h00003DDA: begin
				q			<=			16'hF65F;
		end
		32'h00003DDC: begin
				q			<=			16'h8793;
		end
		32'h00003DDE: begin
				q			<=			16'h004A;
		end
		32'h00003DE0: begin
				q			<=			16'h2623;
		end
		32'h00003DE2: begin
				q			<=			16'h00F1;
		end
		32'h00003DE4: begin
				q			<=			16'h03A3;
		end
		32'h00003DE6: begin
				q			<=			16'h0A01;
		end
		32'h00003DE8: begin
				q			<=			16'h0793;
		end
		32'h00003DEA: begin
				q			<=			16'hFFF0;
		end
		32'h00003DEC: begin
				q			<=			16'h2023;
		end
		32'h00003DEE: begin
				q			<=			16'h0311;
		end
		32'h00003DF0: begin
				q			<=			16'hA483;
		end
		32'h00003DF2: begin
				q			<=			16'h000A;
		end
		32'h00003DF4: begin
				q			<=			16'h0663;
		end
		32'h00003DF6: begin
				q			<=			16'h02FB;
		end
		32'h00003DF8: begin
				q			<=			16'h0613;
		end
		32'h00003DFA: begin
				q			<=			16'h000B;
		end
		32'h00003DFC: begin
				q			<=			16'h0593;
		end
		32'h00003DFE: begin
				q			<=			16'h0000;
		end
		32'h00003E00: begin
				q			<=			16'h8513;
		end
		32'h00003E02: begin
				q			<=			16'h0004;
		end
		32'h00003E04: begin
				q			<=			16'h30EF;
		end
		32'h00003E06: begin
				q			<=			16'h4550;
		end
		32'h00003E08: begin
				q			<=			16'h2223;
		end
		32'h00003E0A: begin
				q			<=			16'h00A1;
		end
		32'h00003E0C: begin
				q			<=			16'h2883;
		end
		32'h00003E0E: begin
				q			<=			16'h0201;
		end
		32'h00003E10: begin
				q			<=			16'h0E63;
		end
		32'h00003E12: begin
				q			<=			16'hE005;
		end
		32'h00003E14: begin
				q			<=			16'h0B33;
		end
		32'h00003E16: begin
				q			<=			16'h4095;
		end
		32'h00003E18: begin
				q			<=			16'h2223;
		end
		32'h00003E1A: begin
				q			<=			16'h0001;
		end
		32'h00003E1C: begin
				q			<=			16'hF06F;
		end
		32'h00003E1E: begin
				q			<=			16'hE10F;
		end
		32'h00003E20: begin
				q			<=			16'h8513;
		end
		32'h00003E22: begin
				q			<=			16'h0004;
		end
		32'h00003E24: begin
				q			<=			16'hF0EF;
		end
		32'h00003E26: begin
				q			<=			16'h808F;
		end
		32'h00003E28: begin
				q			<=			16'h2883;
		end
		32'h00003E2A: begin
				q			<=			16'h0201;
		end
		32'h00003E2C: begin
				q			<=			16'h0B13;
		end
		32'h00003E2E: begin
				q			<=			16'h0005;
		end
		32'h00003E30: begin
				q			<=			16'h2223;
		end
		32'h00003E32: begin
				q			<=			16'h0001;
		end
		32'h00003E34: begin
				q			<=			16'h0D93;
		end
		32'h00003E36: begin
				q			<=			16'h0000;
		end
		32'h00003E38: begin
				q			<=			16'h0C13;
		end
		32'h00003E3A: begin
				q			<=			16'h0000;
		end
		32'h00003E3C: begin
				q			<=			16'h0B93;
		end
		32'h00003E3E: begin
				q			<=			16'h0000;
		end
		32'h00003E40: begin
				q			<=			16'h0C93;
		end
		32'h00003E42: begin
				q			<=			16'h0000;
		end
		32'h00003E44: begin
				q			<=			16'h2023;
		end
		32'h00003E46: begin
				q			<=			16'h03B1;
		end
		32'h00003E48: begin
				q			<=			16'hD463;
		end
		32'h00003E4A: begin
				q			<=			16'h016D;
		end
		32'h00003E4C: begin
				q			<=			16'h2023;
		end
		32'h00003E4E: begin
				q			<=			16'h0361;
		end
		32'h00003E50: begin
				q			<=			16'h4703;
		end
		32'h00003E52: begin
				q			<=			16'h0A71;
		end
		32'h00003E54: begin
				q			<=			16'h0863;
		end
		32'h00003E56: begin
				q			<=			16'h0007;
		end
		32'h00003E58: begin
				q			<=			16'h2783;
		end
		32'h00003E5A: begin
				q			<=			16'h0201;
		end
		32'h00003E5C: begin
				q			<=			16'h8793;
		end
		32'h00003E5E: begin
				q			<=			16'h0017;
		end
		32'h00003E60: begin
				q			<=			16'h2023;
		end
		32'h00003E62: begin
				q			<=			16'h02F1;
		end
		32'h00003E64: begin
				q			<=			16'h7793;
		end
		32'h00003E66: begin
				q			<=			16'h0024;
		end
		32'h00003E68: begin
				q			<=			16'h2C23;
		end
		32'h00003E6A: begin
				q			<=			16'h02F1;
		end
		32'h00003E6C: begin
				q			<=			16'h8863;
		end
		32'h00003E6E: begin
				q			<=			16'h0007;
		end
		32'h00003E70: begin
				q			<=			16'h2783;
		end
		32'h00003E72: begin
				q			<=			16'h0201;
		end
		32'h00003E74: begin
				q			<=			16'h8793;
		end
		32'h00003E76: begin
				q			<=			16'h0027;
		end
		32'h00003E78: begin
				q			<=			16'h2023;
		end
		32'h00003E7A: begin
				q			<=			16'h02F1;
		end
		32'h00003E7C: begin
				q			<=			16'h7A93;
		end
		32'h00003E7E: begin
				q			<=			16'h0844;
		end
		32'h00003E80: begin
				q			<=			16'h9863;
		end
		32'h00003E82: begin
				q			<=			16'h060A;
		end
		32'h00003E84: begin
				q			<=			16'h2783;
		end
		32'h00003E86: begin
				q			<=			16'h01C1;
		end
		32'h00003E88: begin
				q			<=			16'h2703;
		end
		32'h00003E8A: begin
				q			<=			16'h0201;
		end
		32'h00003E8C: begin
				q			<=			16'h8E33;
		end
		32'h00003E8E: begin
				q			<=			16'h40E7;
		end
		32'h00003E90: begin
				q			<=			16'h5063;
		end
		32'h00003E92: begin
				q			<=			16'h07C0;
		end
		32'h00003E94: begin
				q			<=			16'h0F13;
		end
		32'h00003E96: begin
				q			<=			16'h0100;
		end
		32'h00003E98: begin
				q			<=			16'hBE97;
		end
		32'h00003E9A: begin
				q			<=			16'h0000;
		end
		32'h00003E9C: begin
				q			<=			16'h8E93;
		end
		32'h00003E9E: begin
				q			<=			16'h3F4E;
		end
		32'h00003EA0: begin
				q			<=			16'h0F93;
		end
		32'h00003EA2: begin
				q			<=			16'h0070;
		end
		32'h00003EA4: begin
				q			<=			16'h2683;
		end
		32'h00003EA6: begin
				q			<=			16'h0C81;
		end
		32'h00003EA8: begin
				q			<=			16'hA023;
		end
		32'h00003EAA: begin
				q			<=			16'h01D8;
		end
		32'h00003EAC: begin
				q			<=			16'h2703;
		end
		32'h00003EAE: begin
				q			<=			16'h0CC1;
		end
		32'h00003EB0: begin
				q			<=			16'h8693;
		end
		32'h00003EB2: begin
				q			<=			16'h0016;
		end
		32'h00003EB4: begin
				q			<=			16'h8613;
		end
		32'h00003EB6: begin
				q			<=			16'h0088;
		end
		32'h00003EB8: begin
				q			<=			16'h4A63;
		end
		32'h00003EBA: begin
				q			<=			16'h47CF;
		end
		32'h00003EBC: begin
				q			<=			16'h0733;
		end
		32'h00003EBE: begin
				q			<=			16'h00EE;
		end
		32'h00003EC0: begin
				q			<=			16'hA223;
		end
		32'h00003EC2: begin
				q			<=			16'h01C8;
		end
		32'h00003EC4: begin
				q			<=			16'h2623;
		end
		32'h00003EC6: begin
				q			<=			16'h0CE1;
		end
		32'h00003EC8: begin
				q			<=			16'h2423;
		end
		32'h00003ECA: begin
				q			<=			16'h0CD1;
		end
		32'h00003ECC: begin
				q			<=			16'h0713;
		end
		32'h00003ECE: begin
				q			<=			16'h0070;
		end
		32'h00003ED0: begin
				q			<=			16'h0893;
		end
		32'h00003ED2: begin
				q			<=			16'h0006;
		end
		32'h00003ED4: begin
				q			<=			16'h5E63;
		end
		32'h00003ED6: begin
				q			<=			16'h00D7;
		end
		32'h00003ED8: begin
				q			<=			16'h0613;
		end
		32'h00003EDA: begin
				q			<=			16'h0C41;
		end
		32'h00003EDC: begin
				q			<=			16'h8593;
		end
		32'h00003EDE: begin
				q			<=			16'h0009;
		end
		32'h00003EE0: begin
				q			<=			16'h0513;
		end
		32'h00003EE2: begin
				q			<=			16'h0009;
		end
		32'h00003EE4: begin
				q			<=			16'h40EF;
		end
		32'h00003EE6: begin
				q			<=			16'h4790;
		end
		32'h00003EE8: begin
				q			<=			16'h14E3;
		end
		32'h00003EEA: begin
				q			<=			16'h6C05;
		end
		32'h00003EEC: begin
				q			<=			16'h0893;
		end
		32'h00003EEE: begin
				q			<=			16'h0EC1;
		end
		32'h00003EF0: begin
				q			<=			16'h4703;
		end
		32'h00003EF2: begin
				q			<=			16'h0A71;
		end
		32'h00003EF4: begin
				q			<=			16'h0863;
		end
		32'h00003EF6: begin
				q			<=			16'h0407;
		end
		32'h00003EF8: begin
				q			<=			16'h0713;
		end
		32'h00003EFA: begin
				q			<=			16'h0A71;
		end
		32'h00003EFC: begin
				q			<=			16'hA023;
		end
		32'h00003EFE: begin
				q			<=			16'h00E8;
		end
		32'h00003F00: begin
				q			<=			16'h0713;
		end
		32'h00003F02: begin
				q			<=			16'h0010;
		end
		32'h00003F04: begin
				q			<=			16'hA223;
		end
		32'h00003F06: begin
				q			<=			16'h00E8;
		end
		32'h00003F08: begin
				q			<=			16'h2703;
		end
		32'h00003F0A: begin
				q			<=			16'h0CC1;
		end
		32'h00003F0C: begin
				q			<=			16'h0693;
		end
		32'h00003F0E: begin
				q			<=			16'h0070;
		end
		32'h00003F10: begin
				q			<=			16'h8893;
		end
		32'h00003F12: begin
				q			<=			16'h0088;
		end
		32'h00003F14: begin
				q			<=			16'h0713;
		end
		32'h00003F16: begin
				q			<=			16'h0017;
		end
		32'h00003F18: begin
				q			<=			16'h2623;
		end
		32'h00003F1A: begin
				q			<=			16'h0CE1;
		end
		32'h00003F1C: begin
				q			<=			16'h2703;
		end
		32'h00003F1E: begin
				q			<=			16'h0C81;
		end
		32'h00003F20: begin
				q			<=			16'h0713;
		end
		32'h00003F22: begin
				q			<=			16'h0017;
		end
		32'h00003F24: begin
				q			<=			16'h2423;
		end
		32'h00003F26: begin
				q			<=			16'h0CE1;
		end
		32'h00003F28: begin
				q			<=			16'hDE63;
		end
		32'h00003F2A: begin
				q			<=			16'h00E6;
		end
		32'h00003F2C: begin
				q			<=			16'h0613;
		end
		32'h00003F2E: begin
				q			<=			16'h0C41;
		end
		32'h00003F30: begin
				q			<=			16'h8593;
		end
		32'h00003F32: begin
				q			<=			16'h0009;
		end
		32'h00003F34: begin
				q			<=			16'h0513;
		end
		32'h00003F36: begin
				q			<=			16'h0009;
		end
		32'h00003F38: begin
				q			<=			16'h40EF;
		end
		32'h00003F3A: begin
				q			<=			16'h4250;
		end
		32'h00003F3C: begin
				q			<=			16'h1AE3;
		end
		32'h00003F3E: begin
				q			<=			16'h6605;
		end
		32'h00003F40: begin
				q			<=			16'h0893;
		end
		32'h00003F42: begin
				q			<=			16'h0EC1;
		end
		32'h00003F44: begin
				q			<=			16'h2783;
		end
		32'h00003F46: begin
				q			<=			16'h0381;
		end
		32'h00003F48: begin
				q			<=			16'h8863;
		end
		32'h00003F4A: begin
				q			<=			16'h0407;
		end
		32'h00003F4C: begin
				q			<=			16'h0713;
		end
		32'h00003F4E: begin
				q			<=			16'h0A81;
		end
		32'h00003F50: begin
				q			<=			16'hA023;
		end
		32'h00003F52: begin
				q			<=			16'h00E8;
		end
		32'h00003F54: begin
				q			<=			16'h0713;
		end
		32'h00003F56: begin
				q			<=			16'h0020;
		end
		32'h00003F58: begin
				q			<=			16'hA223;
		end
		32'h00003F5A: begin
				q			<=			16'h00E8;
		end
		32'h00003F5C: begin
				q			<=			16'h2703;
		end
		32'h00003F5E: begin
				q			<=			16'h0CC1;
		end
		32'h00003F60: begin
				q			<=			16'h0693;
		end
		32'h00003F62: begin
				q			<=			16'h0070;
		end
		32'h00003F64: begin
				q			<=			16'h8893;
		end
		32'h00003F66: begin
				q			<=			16'h0088;
		end
		32'h00003F68: begin
				q			<=			16'h0713;
		end
		32'h00003F6A: begin
				q			<=			16'h0027;
		end
		32'h00003F6C: begin
				q			<=			16'h2623;
		end
		32'h00003F6E: begin
				q			<=			16'h0CE1;
		end
		32'h00003F70: begin
				q			<=			16'h2703;
		end
		32'h00003F72: begin
				q			<=			16'h0C81;
		end
		32'h00003F74: begin
				q			<=			16'h0713;
		end
		32'h00003F76: begin
				q			<=			16'h0017;
		end
		32'h00003F78: begin
				q			<=			16'h2423;
		end
		32'h00003F7A: begin
				q			<=			16'h0CE1;
		end
		32'h00003F7C: begin
				q			<=			16'hDE63;
		end
		32'h00003F7E: begin
				q			<=			16'h00E6;
		end
		32'h00003F80: begin
				q			<=			16'h0613;
		end
		32'h00003F82: begin
				q			<=			16'h0C41;
		end
		32'h00003F84: begin
				q			<=			16'h8593;
		end
		32'h00003F86: begin
				q			<=			16'h0009;
		end
		32'h00003F88: begin
				q			<=			16'h0513;
		end
		32'h00003F8A: begin
				q			<=			16'h0009;
		end
		32'h00003F8C: begin
				q			<=			16'h40EF;
		end
		32'h00003F8E: begin
				q			<=			16'h3D10;
		end
		32'h00003F90: begin
				q			<=			16'h10E3;
		end
		32'h00003F92: begin
				q			<=			16'h6205;
		end
		32'h00003F94: begin
				q			<=			16'h0893;
		end
		32'h00003F96: begin
				q			<=			16'h0EC1;
		end
		32'h00003F98: begin
				q			<=			16'h0713;
		end
		32'h00003F9A: begin
				q			<=			16'h0800;
		end
		32'h00003F9C: begin
				q			<=			16'h9863;
		end
		32'h00003F9E: begin
				q			<=			16'h06EA;
		end
		32'h00003FA0: begin
				q			<=			16'h2783;
		end
		32'h00003FA2: begin
				q			<=			16'h01C1;
		end
		32'h00003FA4: begin
				q			<=			16'h2703;
		end
		32'h00003FA6: begin
				q			<=			16'h0201;
		end
		32'h00003FA8: begin
				q			<=			16'h8AB3;
		end
		32'h00003FAA: begin
				q			<=			16'h40E7;
		end
		32'h00003FAC: begin
				q			<=			16'h5063;
		end
		32'h00003FAE: begin
				q			<=			16'h0750;
		end
		32'h00003FB0: begin
				q			<=			16'h0E13;
		end
		32'h00003FB2: begin
				q			<=			16'h0100;
		end
		32'h00003FB4: begin
				q			<=			16'hB797;
		end
		32'h00003FB6: begin
				q			<=			16'h0000;
		end
		32'h00003FB8: begin
				q			<=			16'h8793;
		end
		32'h00003FBA: begin
				q			<=			16'h2E87;
		end
		32'h00003FBC: begin
				q			<=			16'h0E93;
		end
		32'h00003FBE: begin
				q			<=			16'h0070;
		end
		32'h00003FC0: begin
				q			<=			16'h2683;
		end
		32'h00003FC2: begin
				q			<=			16'h0C81;
		end
		32'h00003FC4: begin
				q			<=			16'hA023;
		end
		32'h00003FC6: begin
				q			<=			16'h00F8;
		end
		32'h00003FC8: begin
				q			<=			16'h2703;
		end
		32'h00003FCA: begin
				q			<=			16'h0CC1;
		end
		32'h00003FCC: begin
				q			<=			16'h8693;
		end
		32'h00003FCE: begin
				q			<=			16'h0016;
		end
		32'h00003FD0: begin
				q			<=			16'h8613;
		end
		32'h00003FD2: begin
				q			<=			16'h0088;
		end
		32'h00003FD4: begin
				q			<=			16'h4863;
		end
		32'h00003FD6: begin
				q			<=			16'h3B5E;
		end
		32'h00003FD8: begin
				q			<=			16'h8733;
		end
		32'h00003FDA: begin
				q			<=			16'h00EA;
		end
		32'h00003FDC: begin
				q			<=			16'hA223;
		end
		32'h00003FDE: begin
				q			<=			16'h0158;
		end
		32'h00003FE0: begin
				q			<=			16'h2623;
		end
		32'h00003FE2: begin
				q			<=			16'h0CE1;
		end
		32'h00003FE4: begin
				q			<=			16'h2423;
		end
		32'h00003FE6: begin
				q			<=			16'h0CD1;
		end
		32'h00003FE8: begin
				q			<=			16'h0713;
		end
		32'h00003FEA: begin
				q			<=			16'h0070;
		end
		32'h00003FEC: begin
				q			<=			16'h0893;
		end
		32'h00003FEE: begin
				q			<=			16'h0006;
		end
		32'h00003FF0: begin
				q			<=			16'h5E63;
		end
		32'h00003FF2: begin
				q			<=			16'h00D7;
		end
		32'h00003FF4: begin
				q			<=			16'h0613;
		end
		32'h00003FF6: begin
				q			<=			16'h0C41;
		end
		32'h00003FF8: begin
				q			<=			16'h8593;
		end
		32'h00003FFA: begin
				q			<=			16'h0009;
		end
		32'h00003FFC: begin
				q			<=			16'h0513;
		end
		32'h00003FFE: begin
				q			<=			16'h0009;
		end
		32'h00004000: begin
				q			<=			16'h40EF;
		end
		32'h00004002: begin
				q			<=			16'h35D0;
		end
		32'h00004004: begin
				q			<=			16'h16E3;
		end
		32'h00004006: begin
				q			<=			16'h5A05;
		end
		32'h00004008: begin
				q			<=			16'h0893;
		end
		32'h0000400A: begin
				q			<=			16'h0EC1;
		end
		32'h0000400C: begin
				q			<=			16'h8AB3;
		end
		32'h0000400E: begin
				q			<=			16'h416D;
		end
		32'h00004010: begin
				q			<=			16'h5063;
		end
		32'h00004012: begin
				q			<=			16'h0750;
		end
		32'h00004014: begin
				q			<=			16'h0813;
		end
		32'h00004016: begin
				q			<=			16'h0100;
		end
		32'h00004018: begin
				q			<=			16'hBD97;
		end
		32'h0000401A: begin
				q			<=			16'h0000;
		end
		32'h0000401C: begin
				q			<=			16'h8D93;
		end
		32'h0000401E: begin
				q			<=			16'h284D;
		end
		32'h00004020: begin
				q			<=			16'h0E13;
		end
		32'h00004022: begin
				q			<=			16'h0070;
		end
		32'h00004024: begin
				q			<=			16'h2703;
		end
		32'h00004026: begin
				q			<=			16'h0C81;
		end
		32'h00004028: begin
				q			<=			16'hA023;
		end
		32'h0000402A: begin
				q			<=			16'h01B8;
		end
		32'h0000402C: begin
				q			<=			16'h2683;
		end
		32'h0000402E: begin
				q			<=			16'h0CC1;
		end
		32'h00004030: begin
				q			<=			16'h0713;
		end
		32'h00004032: begin
				q			<=			16'h0017;
		end
		32'h00004034: begin
				q			<=			16'h8613;
		end
		32'h00004036: begin
				q			<=			16'h0088;
		end
		32'h00004038: begin
				q			<=			16'h4E63;
		end
		32'h0000403A: begin
				q			<=			16'h3958;
		end
		32'h0000403C: begin
				q			<=			16'hA223;
		end
		32'h0000403E: begin
				q			<=			16'h0158;
		end
		32'h00004040: begin
				q			<=			16'h8AB3;
		end
		32'h00004042: begin
				q			<=			16'h00DA;
		end
		32'h00004044: begin
				q			<=			16'h2623;
		end
		32'h00004046: begin
				q			<=			16'h0D51;
		end
		32'h00004048: begin
				q			<=			16'h2423;
		end
		32'h0000404A: begin
				q			<=			16'h0CE1;
		end
		32'h0000404C: begin
				q			<=			16'h0693;
		end
		32'h0000404E: begin
				q			<=			16'h0070;
		end
		32'h00004050: begin
				q			<=			16'h0893;
		end
		32'h00004052: begin
				q			<=			16'h0006;
		end
		32'h00004054: begin
				q			<=			16'hDE63;
		end
		32'h00004056: begin
				q			<=			16'h00E6;
		end
		32'h00004058: begin
				q			<=			16'h0613;
		end
		32'h0000405A: begin
				q			<=			16'h0C41;
		end
		32'h0000405C: begin
				q			<=			16'h8593;
		end
		32'h0000405E: begin
				q			<=			16'h0009;
		end
		32'h00004060: begin
				q			<=			16'h0513;
		end
		32'h00004062: begin
				q			<=			16'h0009;
		end
		32'h00004064: begin
				q			<=			16'h40EF;
		end
		32'h00004066: begin
				q			<=			16'h2F90;
		end
		32'h00004068: begin
				q			<=			16'h14E3;
		end
		32'h0000406A: begin
				q			<=			16'h5405;
		end
		32'h0000406C: begin
				q			<=			16'h0893;
		end
		32'h0000406E: begin
				q			<=			16'h0EC1;
		end
		32'h00004070: begin
				q			<=			16'h7713;
		end
		32'h00004072: begin
				q			<=			16'h1004;
		end
		32'h00004074: begin
				q			<=			16'h2D83;
		end
		32'h00004076: begin
				q			<=			16'h0CC1;
		end
		32'h00004078: begin
				q			<=			16'h1263;
		end
		32'h0000407A: begin
				q			<=			16'h3A07;
		end
		32'h0000407C: begin
				q			<=			16'h0333;
		end
		32'h0000407E: begin
				q			<=			16'h01BB;
		end
		32'h00004080: begin
				q			<=			16'hA023;
		end
		32'h00004082: begin
				q			<=			16'h0098;
		end
		32'h00004084: begin
				q			<=			16'hA223;
		end
		32'h00004086: begin
				q			<=			16'h0168;
		end
		32'h00004088: begin
				q			<=			16'h2623;
		end
		32'h0000408A: begin
				q			<=			16'h0C61;
		end
		32'h0000408C: begin
				q			<=			16'h2783;
		end
		32'h0000408E: begin
				q			<=			16'h0C81;
		end
		32'h00004090: begin
				q			<=			16'h0713;
		end
		32'h00004092: begin
				q			<=			16'h0070;
		end
		32'h00004094: begin
				q			<=			16'h8893;
		end
		32'h00004096: begin
				q			<=			16'h0088;
		end
		32'h00004098: begin
				q			<=			16'h8793;
		end
		32'h0000409A: begin
				q			<=			16'h0017;
		end
		32'h0000409C: begin
				q			<=			16'h2423;
		end
		32'h0000409E: begin
				q			<=			16'h0CF1;
		end
		32'h000040A0: begin
				q			<=			16'h5263;
		end
		32'h000040A2: begin
				q			<=			16'h4CF7;
		end
		32'h000040A4: begin
				q			<=			16'h0613;
		end
		32'h000040A6: begin
				q			<=			16'h0C41;
		end
		32'h000040A8: begin
				q			<=			16'h8593;
		end
		32'h000040AA: begin
				q			<=			16'h0009;
		end
		32'h000040AC: begin
				q			<=			16'h0513;
		end
		32'h000040AE: begin
				q			<=			16'h0009;
		end
		32'h000040B0: begin
				q			<=			16'h40EF;
		end
		32'h000040B2: begin
				q			<=			16'h2AD0;
		end
		32'h000040B4: begin
				q			<=			16'h1EE3;
		end
		32'h000040B6: begin
				q			<=			16'h4E05;
		end
		32'h000040B8: begin
				q			<=			16'h0893;
		end
		32'h000040BA: begin
				q			<=			16'h0EC1;
		end
		32'h000040BC: begin
				q			<=			16'h006F;
		end
		32'h000040BE: begin
				q			<=			16'h4A80;
		end
		32'h000040C0: begin
				q			<=			16'h6413;
		end
		32'h000040C2: begin
				q			<=			16'h0104;
		end
		32'h000040C4: begin
				q			<=			16'h7793;
		end
		32'h000040C6: begin
				q			<=			16'h0204;
		end
		32'h000040C8: begin
				q			<=			16'h8263;
		end
		32'h000040CA: begin
				q			<=			16'h0207;
		end
		32'h000040CC: begin
				q			<=			16'h8A93;
		end
		32'h000040CE: begin
				q			<=			16'h007A;
		end
		32'h000040D0: begin
				q			<=			16'hFA93;
		end
		32'h000040D2: begin
				q			<=			16'hFF8A;
		end
		32'h000040D4: begin
				q			<=			16'hAC03;
		end
		32'h000040D6: begin
				q			<=			16'h000A;
		end
		32'h000040D8: begin
				q			<=			16'hAC83;
		end
		32'h000040DA: begin
				q			<=			16'h004A;
		end
		32'h000040DC: begin
				q			<=			16'h8793;
		end
		32'h000040DE: begin
				q			<=			16'h008A;
		end
		32'h000040E0: begin
				q			<=			16'h2623;
		end
		32'h000040E2: begin
				q			<=			16'h00F1;
		end
		32'h000040E4: begin
				q			<=			16'h0793;
		end
		32'h000040E6: begin
				q			<=			16'h0010;
		end
		32'h000040E8: begin
				q			<=			16'hF06F;
		end
		32'h000040EA: begin
				q			<=			16'hC55F;
		end
		32'h000040EC: begin
				q			<=			16'h8793;
		end
		32'h000040EE: begin
				q			<=			16'h004A;
		end
		32'h000040F0: begin
				q			<=			16'h2623;
		end
		32'h000040F2: begin
				q			<=			16'h00F1;
		end
		32'h000040F4: begin
				q			<=			16'h7793;
		end
		32'h000040F6: begin
				q			<=			16'h0104;
		end
		32'h000040F8: begin
				q			<=			16'h8663;
		end
		32'h000040FA: begin
				q			<=			16'h0007;
		end
		32'h000040FC: begin
				q			<=			16'hAC03;
		end
		32'h000040FE: begin
				q			<=			16'h000A;
		end
		32'h00004100: begin
				q			<=			16'h006F;
		end
		32'h00004102: begin
				q			<=			16'h0100;
		end
		32'h00004104: begin
				q			<=			16'h7793;
		end
		32'h00004106: begin
				q			<=			16'h0404;
		end
		32'h00004108: begin
				q			<=			16'h8863;
		end
		32'h0000410A: begin
				q			<=			16'h0007;
		end
		32'h0000410C: begin
				q			<=			16'hDC03;
		end
		32'h0000410E: begin
				q			<=			16'h000A;
		end
		32'h00004110: begin
				q			<=			16'h0C93;
		end
		32'h00004112: begin
				q			<=			16'h0000;
		end
		32'h00004114: begin
				q			<=			16'hF06F;
		end
		32'h00004116: begin
				q			<=			16'hFD1F;
		end
		32'h00004118: begin
				q			<=			16'h7793;
		end
		32'h0000411A: begin
				q			<=			16'h2004;
		end
		32'h0000411C: begin
				q			<=			16'h80E3;
		end
		32'h0000411E: begin
				q			<=			16'hFE07;
		end
		32'h00004120: begin
				q			<=			16'hCC03;
		end
		32'h00004122: begin
				q			<=			16'h000A;
		end
		32'h00004124: begin
				q			<=			16'hF06F;
		end
		32'h00004126: begin
				q			<=			16'hFEDF;
		end
		32'h00004128: begin
				q			<=			16'hC797;
		end
		32'h0000412A: begin
				q			<=			16'h0000;
		end
		32'h0000412C: begin
				q			<=			16'h8793;
		end
		32'h0000412E: begin
				q			<=			16'hC5C7;
		end
		32'h00004130: begin
				q			<=			16'hE06F;
		end
		32'h00004132: begin
				q			<=			16'hF75F;
		end
		32'h00004134: begin
				q			<=			16'h8793;
		end
		32'h00004136: begin
				q			<=			16'h004A;
		end
		32'h00004138: begin
				q			<=			16'h2623;
		end
		32'h0000413A: begin
				q			<=			16'h00F1;
		end
		32'h0000413C: begin
				q			<=			16'h7793;
		end
		32'h0000413E: begin
				q			<=			16'h0104;
		end
		32'h00004140: begin
				q			<=			16'h8663;
		end
		32'h00004142: begin
				q			<=			16'h0007;
		end
		32'h00004144: begin
				q			<=			16'hAC03;
		end
		32'h00004146: begin
				q			<=			16'h000A;
		end
		32'h00004148: begin
				q			<=			16'h006F;
		end
		32'h0000414A: begin
				q			<=			16'h0100;
		end
		32'h0000414C: begin
				q			<=			16'h7793;
		end
		32'h0000414E: begin
				q			<=			16'h0404;
		end
		32'h00004150: begin
				q			<=			16'h8863;
		end
		32'h00004152: begin
				q			<=			16'h0007;
		end
		32'h00004154: begin
				q			<=			16'hDC03;
		end
		32'h00004156: begin
				q			<=			16'h000A;
		end
		32'h00004158: begin
				q			<=			16'h0C93;
		end
		32'h0000415A: begin
				q			<=			16'h0000;
		end
		32'h0000415C: begin
				q			<=			16'hE06F;
		end
		32'h0000415E: begin
				q			<=			16'hF71F;
		end
		32'h00004160: begin
				q			<=			16'h7793;
		end
		32'h00004162: begin
				q			<=			16'h2004;
		end
		32'h00004164: begin
				q			<=			16'h80E3;
		end
		32'h00004166: begin
				q			<=			16'hFE07;
		end
		32'h00004168: begin
				q			<=			16'hCC03;
		end
		32'h0000416A: begin
				q			<=			16'h000A;
		end
		32'h0000416C: begin
				q			<=			16'hF06F;
		end
		32'h0000416E: begin
				q			<=			16'hFEDF;
		end
		32'h00004170: begin
				q			<=			16'h0713;
		end
		32'h00004172: begin
				q			<=			16'h0004;
		end
		32'h00004174: begin
				q			<=			16'h0793;
		end
		32'h00004176: begin
				q			<=			16'h0010;
		end
		32'h00004178: begin
				q			<=			16'hF06F;
		end
		32'h0000417A: begin
				q			<=			16'hBD5F;
		end
		32'h0000417C: begin
				q			<=			16'h0713;
		end
		32'h0000417E: begin
				q			<=			16'h0010;
		end
		32'h00004180: begin
				q			<=			16'h8463;
		end
		32'h00004182: begin
				q			<=			16'h98E7;
		end
		32'h00004184: begin
				q			<=			16'h0713;
		end
		32'h00004186: begin
				q			<=			16'h0020;
		end
		32'h00004188: begin
				q			<=			16'h8E63;
		end
		32'h0000418A: begin
				q			<=			16'h12E7;
		end
		32'h0000418C: begin
				q			<=			16'h0793;
		end
		32'h0000418E: begin
				q			<=			16'h1901;
		end
		32'h00004190: begin
				q			<=			16'h9693;
		end
		32'h00004192: begin
				q			<=			16'h01DC;
		end
		32'h00004194: begin
				q			<=			16'h7713;
		end
		32'h00004196: begin
				q			<=			16'h007C;
		end
		32'h00004198: begin
				q			<=			16'h5C13;
		end
		32'h0000419A: begin
				q			<=			16'h003C;
		end
		32'h0000419C: begin
				q			<=			16'h0713;
		end
		32'h0000419E: begin
				q			<=			16'h0307;
		end
		32'h000041A0: begin
				q			<=			16'hEC33;
		end
		32'h000041A2: begin
				q			<=			16'h0186;
		end
		32'h000041A4: begin
				q			<=			16'hDC93;
		end
		32'h000041A6: begin
				q			<=			16'h003C;
		end
		32'h000041A8: begin
				q			<=			16'h8FA3;
		end
		32'h000041AA: begin
				q			<=			16'hFEE7;
		end
		32'h000041AC: begin
				q			<=			16'h66B3;
		end
		32'h000041AE: begin
				q			<=			16'h019C;
		end
		32'h000041B0: begin
				q			<=			16'h8493;
		end
		32'h000041B2: begin
				q			<=			16'hFFF7;
		end
		32'h000041B4: begin
				q			<=			16'h9E63;
		end
		32'h000041B6: begin
				q			<=			16'h0206;
		end
		32'h000041B8: begin
				q			<=			16'h7693;
		end
		32'h000041BA: begin
				q			<=			16'h0014;
		end
		32'h000041BC: begin
				q			<=			16'h8A63;
		end
		32'h000041BE: begin
				q			<=			16'h0006;
		end
		32'h000041C0: begin
				q			<=			16'h0693;
		end
		32'h000041C2: begin
				q			<=			16'h0300;
		end
		32'h000041C4: begin
				q			<=			16'h0663;
		end
		32'h000041C6: begin
				q			<=			16'h00D7;
		end
		32'h000041C8: begin
				q			<=			16'h8FA3;
		end
		32'h000041CA: begin
				q			<=			16'hFED4;
		end
		32'h000041CC: begin
				q			<=			16'h8493;
		end
		32'h000041CE: begin
				q			<=			16'hFFE7;
		end
		32'h000041D0: begin
				q			<=			16'h0793;
		end
		32'h000041D2: begin
				q			<=			16'h1901;
		end
		32'h000041D4: begin
				q			<=			16'h0D93;
		end
		32'h000041D6: begin
				q			<=			16'h000B;
		end
		32'h000041D8: begin
				q			<=			16'h2223;
		end
		32'h000041DA: begin
				q			<=			16'h0001;
		end
		32'h000041DC: begin
				q			<=			16'h8B33;
		end
		32'h000041DE: begin
				q			<=			16'h4097;
		end
		32'h000041E0: begin
				q			<=			16'h0C13;
		end
		32'h000041E2: begin
				q			<=			16'h0000;
		end
		32'h000041E4: begin
				q			<=			16'h0B93;
		end
		32'h000041E6: begin
				q			<=			16'h0000;
		end
		32'h000041E8: begin
				q			<=			16'h0C93;
		end
		32'h000041EA: begin
				q			<=			16'h0000;
		end
		32'h000041EC: begin
				q			<=			16'hF06F;
		end
		32'h000041EE: begin
				q			<=			16'hC59F;
		end
		32'h000041F0: begin
				q			<=			16'h8793;
		end
		32'h000041F2: begin
				q			<=			16'h0004;
		end
		32'h000041F4: begin
				q			<=			16'hF06F;
		end
		32'h000041F6: begin
				q			<=			16'hF9DF;
		end
		32'h000041F8: begin
				q			<=			16'h0A13;
		end
		32'h000041FA: begin
				q			<=			16'h0000;
		end
		32'h000041FC: begin
				q			<=			16'h0D93;
		end
		32'h000041FE: begin
				q			<=			16'h1901;
		end
		32'h00004200: begin
				q			<=			16'h7A93;
		end
		32'h00004202: begin
				q			<=			16'h4004;
		end
		32'h00004204: begin
				q			<=			16'h0B93;
		end
		32'h00004206: begin
				q			<=			16'h0090;
		end
		32'h00004208: begin
				q			<=			16'h0613;
		end
		32'h0000420A: begin
				q			<=			16'h00A0;
		end
		32'h0000420C: begin
				q			<=			16'h0693;
		end
		32'h0000420E: begin
				q			<=			16'h0000;
		end
		32'h00004210: begin
				q			<=			16'h0513;
		end
		32'h00004212: begin
				q			<=			16'h000C;
		end
		32'h00004214: begin
				q			<=			16'h8593;
		end
		32'h00004216: begin
				q			<=			16'h000C;
		end
		32'h00004218: begin
				q			<=			16'h2223;
		end
		32'h0000421A: begin
				q			<=			16'h0111;
		end
		32'h0000421C: begin
				q			<=			16'h60EF;
		end
		32'h0000421E: begin
				q			<=			16'h4C90;
		end
		32'h00004220: begin
				q			<=			16'h0513;
		end
		32'h00004222: begin
				q			<=			16'h0305;
		end
		32'h00004224: begin
				q			<=			16'h8FA3;
		end
		32'h00004226: begin
				q			<=			16'hFEAD;
		end
		32'h00004228: begin
				q			<=			16'h8493;
		end
		32'h0000422A: begin
				q			<=			16'hFFFD;
		end
		32'h0000422C: begin
				q			<=			16'h0A13;
		end
		32'h0000422E: begin
				q			<=			16'h001A;
		end
		32'h00004230: begin
				q			<=			16'h2883;
		end
		32'h00004232: begin
				q			<=			16'h0041;
		end
		32'h00004234: begin
				q			<=			16'h8E63;
		end
		32'h00004236: begin
				q			<=			16'h040A;
		end
		32'h00004238: begin
				q			<=			16'h2783;
		end
		32'h0000423A: begin
				q			<=			16'h0081;
		end
		32'h0000423C: begin
				q			<=			16'hC783;
		end
		32'h0000423E: begin
				q			<=			16'h0007;
		end
		32'h00004240: begin
				q			<=			16'h1863;
		end
		32'h00004242: begin
				q			<=			16'h04FA;
		end
		32'h00004244: begin
				q			<=			16'h0793;
		end
		32'h00004246: begin
				q			<=			16'h0FF0;
		end
		32'h00004248: begin
				q			<=			16'h0463;
		end
		32'h0000424A: begin
				q			<=			16'h04FA;
		end
		32'h0000424C: begin
				q			<=			16'h9463;
		end
		32'h0000424E: begin
				q			<=			16'h000C;
		end
		32'h00004250: begin
				q			<=			16'hF063;
		end
		32'h00004252: begin
				q			<=			16'h058B;
		end
		32'h00004254: begin
				q			<=			16'h2783;
		end
		32'h00004256: begin
				q			<=			16'h0241;
		end
		32'h00004258: begin
				q			<=			16'h2583;
		end
		32'h0000425A: begin
				q			<=			16'h02C1;
		end
		32'h0000425C: begin
				q			<=			16'h2223;
		end
		32'h0000425E: begin
				q			<=			16'h0111;
		end
		32'h00004260: begin
				q			<=			16'h84B3;
		end
		32'h00004262: begin
				q			<=			16'h40F4;
		end
		32'h00004264: begin
				q			<=			16'h8613;
		end
		32'h00004266: begin
				q			<=			16'h0007;
		end
		32'h00004268: begin
				q			<=			16'h8513;
		end
		32'h0000426A: begin
				q			<=			16'h0004;
		end
		32'h0000426C: begin
				q			<=			16'hE0EF;
		end
		32'h0000426E: begin
				q			<=			16'hC21F;
		end
		32'h00004270: begin
				q			<=			16'h2783;
		end
		32'h00004272: begin
				q			<=			16'h0081;
		end
		32'h00004274: begin
				q			<=			16'h0A13;
		end
		32'h00004276: begin
				q			<=			16'h0000;
		end
		32'h00004278: begin
				q			<=			16'h2883;
		end
		32'h0000427A: begin
				q			<=			16'h0041;
		end
		32'h0000427C: begin
				q			<=			16'hC783;
		end
		32'h0000427E: begin
				q			<=			16'h0017;
		end
		32'h00004280: begin
				q			<=			16'h8863;
		end
		32'h00004282: begin
				q			<=			16'h0007;
		end
		32'h00004284: begin
				q			<=			16'h2783;
		end
		32'h00004286: begin
				q			<=			16'h0081;
		end
		32'h00004288: begin
				q			<=			16'h8793;
		end
		32'h0000428A: begin
				q			<=			16'h0017;
		end
		32'h0000428C: begin
				q			<=			16'h2423;
		end
		32'h0000428E: begin
				q			<=			16'h00F1;
		end
		32'h00004290: begin
				q			<=			16'h0513;
		end
		32'h00004292: begin
				q			<=			16'h000C;
		end
		32'h00004294: begin
				q			<=			16'h8593;
		end
		32'h00004296: begin
				q			<=			16'h000C;
		end
		32'h00004298: begin
				q			<=			16'h0613;
		end
		32'h0000429A: begin
				q			<=			16'h00A0;
		end
		32'h0000429C: begin
				q			<=			16'h0693;
		end
		32'h0000429E: begin
				q			<=			16'h0000;
		end
		32'h000042A0: begin
				q			<=			16'h2223;
		end
		32'h000042A2: begin
				q			<=			16'h0111;
		end
		32'h000042A4: begin
				q			<=			16'h60EF;
		end
		32'h000042A6: begin
				q			<=			16'h0090;
		end
		32'h000042A8: begin
				q			<=			16'h8C93;
		end
		32'h000042AA: begin
				q			<=			16'h0005;
		end
		32'h000042AC: begin
				q			<=			16'hE5B3;
		end
		32'h000042AE: begin
				q			<=			16'h00A5;
		end
		32'h000042B0: begin
				q			<=			16'h0C13;
		end
		32'h000042B2: begin
				q			<=			16'h0005;
		end
		32'h000042B4: begin
				q			<=			16'h2883;
		end
		32'h000042B6: begin
				q			<=			16'h0041;
		end
		32'h000042B8: begin
				q			<=			16'h8CE3;
		end
		32'h000042BA: begin
				q			<=			16'hF005;
		end
		32'h000042BC: begin
				q			<=			16'h8D93;
		end
		32'h000042BE: begin
				q			<=			16'h0004;
		end
		32'h000042C0: begin
				q			<=			16'hF06F;
		end
		32'h000042C2: begin
				q			<=			16'hF49F;
		end
		32'h000042C4: begin
				q			<=			16'h0493;
		end
		32'h000042C6: begin
				q			<=			16'h1901;
		end
		32'h000042C8: begin
				q			<=			16'h2703;
		end
		32'h000042CA: begin
				q			<=			16'h0341;
		end
		32'h000042CC: begin
				q			<=			16'h7793;
		end
		32'h000042CE: begin
				q			<=			16'h00FC;
		end
		32'h000042D0: begin
				q			<=			16'h8493;
		end
		32'h000042D2: begin
				q			<=			16'hFFF4;
		end
		32'h000042D4: begin
				q			<=			16'h07B3;
		end
		32'h000042D6: begin
				q			<=			16'h00F7;
		end
		32'h000042D8: begin
				q			<=			16'hC783;
		end
		32'h000042DA: begin
				q			<=			16'h0007;
		end
		32'h000042DC: begin
				q			<=			16'h5C13;
		end
		32'h000042DE: begin
				q			<=			16'h004C;
		end
		32'h000042E0: begin
				q			<=			16'h8023;
		end
		32'h000042E2: begin
				q			<=			16'h00F4;
		end
		32'h000042E4: begin
				q			<=			16'h9793;
		end
		32'h000042E6: begin
				q			<=			16'h01CC;
		end
		32'h000042E8: begin
				q			<=			16'hEC33;
		end
		32'h000042EA: begin
				q			<=			16'h0187;
		end
		32'h000042EC: begin
				q			<=			16'hDC93;
		end
		32'h000042EE: begin
				q			<=			16'h004C;
		end
		32'h000042F0: begin
				q			<=			16'h67B3;
		end
		32'h000042F2: begin
				q			<=			16'h019C;
		end
		32'h000042F4: begin
				q			<=			16'h9AE3;
		end
		32'h000042F6: begin
				q			<=			16'hFC07;
		end
		32'h000042F8: begin
				q			<=			16'hF06F;
		end
		32'h000042FA: begin
				q			<=			16'hED9F;
		end
		32'h000042FC: begin
				q			<=			16'h0493;
		end
		32'h000042FE: begin
				q			<=			16'h1901;
		end
		32'h00004300: begin
				q			<=			16'h98E3;
		end
		32'h00004302: begin
				q			<=			16'hEC07;
		end
		32'h00004304: begin
				q			<=			16'h7713;
		end
		32'h00004306: begin
				q			<=			16'h0017;
		end
		32'h00004308: begin
				q			<=			16'h04E3;
		end
		32'h0000430A: begin
				q			<=			16'hEC07;
		end
		32'h0000430C: begin
				q			<=			16'h0793;
		end
		32'h0000430E: begin
				q			<=			16'h0300;
		end
		32'h00004310: begin
				q			<=			16'h07A3;
		end
		32'h00004312: begin
				q			<=			16'h18F1;
		end
		32'h00004314: begin
				q			<=			16'hF06F;
		end
		32'h00004316: begin
				q			<=			16'h808F;
		end
		32'h00004318: begin
				q			<=			16'h02E3;
		end
		32'h0000431A: begin
				q			<=			16'h300D;
		end
		32'h0000431C: begin
				q			<=			16'h0623;
		end
		32'h0000431E: begin
				q			<=			16'h13A1;
		end
		32'h00004320: begin
				q			<=			16'h03A3;
		end
		32'h00004322: begin
				q			<=			16'h0A01;
		end
		32'h00004324: begin
				q			<=			16'h2623;
		end
		32'h00004326: begin
				q			<=			16'h0151;
		end
		32'h00004328: begin
				q			<=			16'hE06F;
		end
		32'h0000432A: begin
				q			<=			16'hF79F;
		end
		32'h0000432C: begin
				q			<=			16'h0713;
		end
		32'h0000432E: begin
				q			<=			16'h0107;
		end
		32'h00004330: begin
				q			<=			16'hA223;
		end
		32'h00004332: begin
				q			<=			16'h01E8;
		end
		32'h00004334: begin
				q			<=			16'h2623;
		end
		32'h00004336: begin
				q			<=			16'h0CE1;
		end
		32'h00004338: begin
				q			<=			16'h2423;
		end
		32'h0000433A: begin
				q			<=			16'h0CD1;
		end
		32'h0000433C: begin
				q			<=			16'hDE63;
		end
		32'h0000433E: begin
				q			<=			16'h02DF;
		end
		32'h00004340: begin
				q			<=			16'h0613;
		end
		32'h00004342: begin
				q			<=			16'h0C41;
		end
		32'h00004344: begin
				q			<=			16'h8593;
		end
		32'h00004346: begin
				q			<=			16'h0009;
		end
		32'h00004348: begin
				q			<=			16'h0513;
		end
		32'h0000434A: begin
				q			<=			16'h0009;
		end
		32'h0000434C: begin
				q			<=			16'h2423;
		end
		32'h0000434E: begin
				q			<=			16'h05F1;
		end
		32'h00004350: begin
				q			<=			16'h2223;
		end
		32'h00004352: begin
				q			<=			16'h05D1;
		end
		32'h00004354: begin
				q			<=			16'h2023;
		end
		32'h00004356: begin
				q			<=			16'h05E1;
		end
		32'h00004358: begin
				q			<=			16'h2E23;
		end
		32'h0000435A: begin
				q			<=			16'h03C1;
		end
		32'h0000435C: begin
				q			<=			16'h40EF;
		end
		32'h0000435E: begin
				q			<=			16'h0010;
		end
		32'h00004360: begin
				q			<=			16'h18E3;
		end
		32'h00004362: begin
				q			<=			16'h2405;
		end
		32'h00004364: begin
				q			<=			16'h2F83;
		end
		32'h00004366: begin
				q			<=			16'h0481;
		end
		32'h00004368: begin
				q			<=			16'h2E83;
		end
		32'h0000436A: begin
				q			<=			16'h0441;
		end
		32'h0000436C: begin
				q			<=			16'h2F03;
		end
		32'h0000436E: begin
				q			<=			16'h0401;
		end
		32'h00004370: begin
				q			<=			16'h2E03;
		end
		32'h00004372: begin
				q			<=			16'h03C1;
		end
		32'h00004374: begin
				q			<=			16'h0613;
		end
		32'h00004376: begin
				q			<=			16'h0EC1;
		end
		32'h00004378: begin
				q			<=			16'h0E13;
		end
		32'h0000437A: begin
				q			<=			16'hFF0E;
		end
		32'h0000437C: begin
				q			<=			16'h0893;
		end
		32'h0000437E: begin
				q			<=			16'h0006;
		end
		32'h00004380: begin
				q			<=			16'hF06F;
		end
		32'h00004382: begin
				q			<=			16'hB25F;
		end
		32'h00004384: begin
				q			<=			16'h0713;
		end
		32'h00004386: begin
				q			<=			16'h0107;
		end
		32'h00004388: begin
				q			<=			16'hA223;
		end
		32'h0000438A: begin
				q			<=			16'h01C8;
		end
		32'h0000438C: begin
				q			<=			16'h2623;
		end
		32'h0000438E: begin
				q			<=			16'h0CE1;
		end
		32'h00004390: begin
				q			<=			16'h2423;
		end
		32'h00004392: begin
				q			<=			16'h0CD1;
		end
		32'h00004394: begin
				q			<=			16'hDA63;
		end
		32'h00004396: begin
				q			<=			16'h02DE;
		end
		32'h00004398: begin
				q			<=			16'h0613;
		end
		32'h0000439A: begin
				q			<=			16'h0C41;
		end
		32'h0000439C: begin
				q			<=			16'h8593;
		end
		32'h0000439E: begin
				q			<=			16'h0009;
		end
		32'h000043A0: begin
				q			<=			16'h0513;
		end
		32'h000043A2: begin
				q			<=			16'h0009;
		end
		32'h000043A4: begin
				q			<=			16'h2023;
		end
		32'h000043A6: begin
				q			<=			16'h05D1;
		end
		32'h000043A8: begin
				q			<=			16'h2E23;
		end
		32'h000043AA: begin
				q			<=			16'h02F1;
		end
		32'h000043AC: begin
				q			<=			16'h2C23;
		end
		32'h000043AE: begin
				q			<=			16'h03C1;
		end
		32'h000043B0: begin
				q			<=			16'h40EF;
		end
		32'h000043B2: begin
				q			<=			16'h7AC0;
		end
		32'h000043B4: begin
				q			<=			16'h1EE3;
		end
		32'h000043B6: begin
				q			<=			16'h1E05;
		end
		32'h000043B8: begin
				q			<=			16'h2E83;
		end
		32'h000043BA: begin
				q			<=			16'h0401;
		end
		32'h000043BC: begin
				q			<=			16'h2783;
		end
		32'h000043BE: begin
				q			<=			16'h03C1;
		end
		32'h000043C0: begin
				q			<=			16'h2E03;
		end
		32'h000043C2: begin
				q			<=			16'h0381;
		end
		32'h000043C4: begin
				q			<=			16'h0613;
		end
		32'h000043C6: begin
				q			<=			16'h0EC1;
		end
		32'h000043C8: begin
				q			<=			16'h8A93;
		end
		32'h000043CA: begin
				q			<=			16'hFF0A;
		end
		32'h000043CC: begin
				q			<=			16'h0893;
		end
		32'h000043CE: begin
				q			<=			16'h0006;
		end
		32'h000043D0: begin
				q			<=			16'hF06F;
		end
		32'h000043D2: begin
				q			<=			16'hBF1F;
		end
		32'h000043D4: begin
				q			<=			16'h8693;
		end
		32'h000043D6: begin
				q			<=			16'h0106;
		end
		32'h000043D8: begin
				q			<=			16'hA223;
		end
		32'h000043DA: begin
				q			<=			16'h0108;
		end
		32'h000043DC: begin
				q			<=			16'h2623;
		end
		32'h000043DE: begin
				q			<=			16'h0CD1;
		end
		32'h000043E0: begin
				q			<=			16'h2423;
		end
		32'h000043E2: begin
				q			<=			16'h0CE1;
		end
		32'h000043E4: begin
				q			<=			16'h5663;
		end
		32'h000043E6: begin
				q			<=			16'h02EE;
		end
		32'h000043E8: begin
				q			<=			16'h0613;
		end
		32'h000043EA: begin
				q			<=			16'h0C41;
		end
		32'h000043EC: begin
				q			<=			16'h8593;
		end
		32'h000043EE: begin
				q			<=			16'h0009;
		end
		32'h000043F0: begin
				q			<=			16'h0513;
		end
		32'h000043F2: begin
				q			<=			16'h0009;
		end
		32'h000043F4: begin
				q			<=			16'h2E23;
		end
		32'h000043F6: begin
				q			<=			16'h03C1;
		end
		32'h000043F8: begin
				q			<=			16'h2C23;
		end
		32'h000043FA: begin
				q			<=			16'h0301;
		end
		32'h000043FC: begin
				q			<=			16'h40EF;
		end
		32'h000043FE: begin
				q			<=			16'h7600;
		end
		32'h00004400: begin
				q			<=			16'h18E3;
		end
		32'h00004402: begin
				q			<=			16'h1A05;
		end
		32'h00004404: begin
				q			<=			16'h2E03;
		end
		32'h00004406: begin
				q			<=			16'h03C1;
		end
		32'h00004408: begin
				q			<=			16'h2803;
		end
		32'h0000440A: begin
				q			<=			16'h0381;
		end
		32'h0000440C: begin
				q			<=			16'h0613;
		end
		32'h0000440E: begin
				q			<=			16'h0EC1;
		end
		32'h00004410: begin
				q			<=			16'h8A93;
		end
		32'h00004412: begin
				q			<=			16'hFF0A;
		end
		32'h00004414: begin
				q			<=			16'h0893;
		end
		32'h00004416: begin
				q			<=			16'h0006;
		end
		32'h00004418: begin
				q			<=			16'hF06F;
		end
		32'h0000441A: begin
				q			<=			16'hC0DF;
		end
		32'h0000441C: begin
				q			<=			16'h0713;
		end
		32'h0000441E: begin
				q			<=			16'h0650;
		end
		32'h00004420: begin
				q			<=			16'h5463;
		end
		32'h00004422: begin
				q			<=			16'h73A7;
		end
		32'h00004424: begin
				q			<=			16'h2703;
		end
		32'h00004426: begin
				q			<=			16'h0D01;
		end
		32'h00004428: begin
				q			<=			16'h0593;
		end
		32'h0000442A: begin
				q			<=			16'h0801;
		end
		32'h0000442C: begin
				q			<=			16'h0513;
		end
		32'h0000442E: begin
				q			<=			16'h0901;
		end
		32'h00004430: begin
				q			<=			16'h2823;
		end
		32'h00004432: begin
				q			<=			16'h08E1;
		end
		32'h00004434: begin
				q			<=			16'h2703;
		end
		32'h00004436: begin
				q			<=			16'h0D41;
		end
		32'h00004438: begin
				q			<=			16'h2C23;
		end
		32'h0000443A: begin
				q			<=			16'h0311;
		end
		32'h0000443C: begin
				q			<=			16'h2023;
		end
		32'h0000443E: begin
				q			<=			16'h0801;
		end
		32'h00004440: begin
				q			<=			16'h2A23;
		end
		32'h00004442: begin
				q			<=			16'h08E1;
		end
		32'h00004444: begin
				q			<=			16'h2703;
		end
		32'h00004446: begin
				q			<=			16'h0D81;
		end
		32'h00004448: begin
				q			<=			16'h2223;
		end
		32'h0000444A: begin
				q			<=			16'h0801;
		end
		32'h0000444C: begin
				q			<=			16'h2423;
		end
		32'h0000444E: begin
				q			<=			16'h0801;
		end
		32'h00004450: begin
				q			<=			16'h2C23;
		end
		32'h00004452: begin
				q			<=			16'h08E1;
		end
		32'h00004454: begin
				q			<=			16'h2703;
		end
		32'h00004456: begin
				q			<=			16'h0DC1;
		end
		32'h00004458: begin
				q			<=			16'h2623;
		end
		32'h0000445A: begin
				q			<=			16'h0801;
		end
		32'h0000445C: begin
				q			<=			16'h2E23;
		end
		32'h0000445E: begin
				q			<=			16'h08E1;
		end
		32'h00004460: begin
				q			<=			16'h70EF;
		end
		32'h00004462: begin
				q			<=			16'h35D0;
		end
		32'h00004464: begin
				q			<=			16'h2883;
		end
		32'h00004466: begin
				q			<=			16'h0381;
		end
		32'h00004468: begin
				q			<=			16'h1463;
		end
		32'h0000446A: begin
				q			<=			16'h1805;
		end
		32'h0000446C: begin
				q			<=			16'hC797;
		end
		32'h0000446E: begin
				q			<=			16'h0000;
		end
		32'h00004470: begin
				q			<=			16'h8793;
		end
		32'h00004472: begin
				q			<=			16'h9407;
		end
		32'h00004474: begin
				q			<=			16'hA023;
		end
		32'h00004476: begin
				q			<=			16'h00F8;
		end
		32'h00004478: begin
				q			<=			16'h0793;
		end
		32'h0000447A: begin
				q			<=			16'h0010;
		end
		32'h0000447C: begin
				q			<=			16'hA223;
		end
		32'h0000447E: begin
				q			<=			16'h00F8;
		end
		32'h00004480: begin
				q			<=			16'h2783;
		end
		32'h00004482: begin
				q			<=			16'h0C81;
		end
		32'h00004484: begin
				q			<=			16'h8D93;
		end
		32'h00004486: begin
				q			<=			16'h001D;
		end
		32'h00004488: begin
				q			<=			16'h2623;
		end
		32'h0000448A: begin
				q			<=			16'h0DB1;
		end
		32'h0000448C: begin
				q			<=			16'h8793;
		end
		32'h0000448E: begin
				q			<=			16'h0017;
		end
		32'h00004490: begin
				q			<=			16'h2423;
		end
		32'h00004492: begin
				q			<=			16'h0CF1;
		end
		32'h00004494: begin
				q			<=			16'h0713;
		end
		32'h00004496: begin
				q			<=			16'h0070;
		end
		32'h00004498: begin
				q			<=			16'h8893;
		end
		32'h0000449A: begin
				q			<=			16'h0088;
		end
		32'h0000449C: begin
				q			<=			16'h5E63;
		end
		32'h0000449E: begin
				q			<=			16'h00F7;
		end
		32'h000044A0: begin
				q			<=			16'h0613;
		end
		32'h000044A2: begin
				q			<=			16'h0C41;
		end
		32'h000044A4: begin
				q			<=			16'h8593;
		end
		32'h000044A6: begin
				q			<=			16'h0009;
		end
		32'h000044A8: begin
				q			<=			16'h0513;
		end
		32'h000044AA: begin
				q			<=			16'h0009;
		end
		32'h000044AC: begin
				q			<=			16'h40EF;
		end
		32'h000044AE: begin
				q			<=			16'h6B00;
		end
		32'h000044B0: begin
				q			<=			16'h10E3;
		end
		32'h000044B2: begin
				q			<=			16'h1005;
		end
		32'h000044B4: begin
				q			<=			16'h0893;
		end
		32'h000044B6: begin
				q			<=			16'h0EC1;
		end
		32'h000044B8: begin
				q			<=			16'h2783;
		end
		32'h000044BA: begin
				q			<=			16'h0AC1;
		end
		32'h000044BC: begin
				q			<=			16'hC663;
		end
		32'h000044BE: begin
				q			<=			16'h0147;
		end
		32'h000044C0: begin
				q			<=			16'h7793;
		end
		32'h000044C2: begin
				q			<=			16'h0014;
		end
		32'h000044C4: begin
				q			<=			16'h8063;
		end
		32'h000044C6: begin
				q			<=			16'h0A07;
		end
		32'h000044C8: begin
				q			<=			16'h2783;
		end
		32'h000044CA: begin
				q			<=			16'h0281;
		end
		32'h000044CC: begin
				q			<=			16'h2703;
		end
		32'h000044CE: begin
				q			<=			16'h0141;
		end
		32'h000044D0: begin
				q			<=			16'h8893;
		end
		32'h000044D2: begin
				q			<=			16'h0088;
		end
		32'h000044D4: begin
				q			<=			16'hAC23;
		end
		32'h000044D6: begin
				q			<=			16'hFEF8;
		end
		32'h000044D8: begin
				q			<=			16'h2783;
		end
		32'h000044DA: begin
				q			<=			16'h0141;
		end
		32'h000044DC: begin
				q			<=			16'hAE23;
		end
		32'h000044DE: begin
				q			<=			16'hFEF8;
		end
		32'h000044E0: begin
				q			<=			16'h2783;
		end
		32'h000044E2: begin
				q			<=			16'h0CC1;
		end
		32'h000044E4: begin
				q			<=			16'h87B3;
		end
		32'h000044E6: begin
				q			<=			16'h00E7;
		end
		32'h000044E8: begin
				q			<=			16'h2623;
		end
		32'h000044EA: begin
				q			<=			16'h0CF1;
		end
		32'h000044EC: begin
				q			<=			16'h2783;
		end
		32'h000044EE: begin
				q			<=			16'h0C81;
		end
		32'h000044F0: begin
				q			<=			16'h0713;
		end
		32'h000044F2: begin
				q			<=			16'h0070;
		end
		32'h000044F4: begin
				q			<=			16'h8793;
		end
		32'h000044F6: begin
				q			<=			16'h0017;
		end
		32'h000044F8: begin
				q			<=			16'h2423;
		end
		32'h000044FA: begin
				q			<=			16'h0CF1;
		end
		32'h000044FC: begin
				q			<=			16'h5E63;
		end
		32'h000044FE: begin
				q			<=			16'h00F7;
		end
		32'h00004500: begin
				q			<=			16'h0613;
		end
		32'h00004502: begin
				q			<=			16'h0C41;
		end
		32'h00004504: begin
				q			<=			16'h8593;
		end
		32'h00004506: begin
				q			<=			16'h0009;
		end
		32'h00004508: begin
				q			<=			16'h0513;
		end
		32'h0000450A: begin
				q			<=			16'h0009;
		end
		32'h0000450C: begin
				q			<=			16'h40EF;
		end
		32'h0000450E: begin
				q			<=			16'h6500;
		end
		32'h00004510: begin
				q			<=			16'h10E3;
		end
		32'h00004512: begin
				q			<=			16'h0A05;
		end
		32'h00004514: begin
				q			<=			16'h0893;
		end
		32'h00004516: begin
				q			<=			16'h0EC1;
		end
		32'h00004518: begin
				q			<=			16'h0493;
		end
		32'h0000451A: begin
				q			<=			16'hFFFA;
		end
		32'h0000451C: begin
				q			<=			16'h5463;
		end
		32'h0000451E: begin
				q			<=			16'h0490;
		end
		32'h00004520: begin
				q			<=			16'h0B93;
		end
		32'h00004522: begin
				q			<=			16'h0100;
		end
		32'h00004524: begin
				q			<=			16'hBA97;
		end
		32'h00004526: begin
				q			<=			16'h0000;
		end
		32'h00004528: begin
				q			<=			16'h8A93;
		end
		32'h0000452A: begin
				q			<=			16'hD78A;
		end
		32'h0000452C: begin
				q			<=			16'h0C13;
		end
		32'h0000452E: begin
				q			<=			16'h0070;
		end
		32'h00004530: begin
				q			<=			16'h2783;
		end
		32'h00004532: begin
				q			<=			16'h0C81;
		end
		32'h00004534: begin
				q			<=			16'hA023;
		end
		32'h00004536: begin
				q			<=			16'h0158;
		end
		32'h00004538: begin
				q			<=			16'h2703;
		end
		32'h0000453A: begin
				q			<=			16'h0CC1;
		end
		32'h0000453C: begin
				q			<=			16'h8793;
		end
		32'h0000453E: begin
				q			<=			16'h0017;
		end
		32'h00004540: begin
				q			<=			16'h8693;
		end
		32'h00004542: begin
				q			<=			16'h0088;
		end
		32'h00004544: begin
				q			<=			16'hCA63;
		end
		32'h00004546: begin
				q			<=			16'h069B;
		end
		32'h00004548: begin
				q			<=			16'hA223;
		end
		32'h0000454A: begin
				q			<=			16'h0098;
		end
		32'h0000454C: begin
				q			<=			16'h84B3;
		end
		32'h0000454E: begin
				q			<=			16'h00E4;
		end
		32'h00004550: begin
				q			<=			16'h2623;
		end
		32'h00004552: begin
				q			<=			16'h0C91;
		end
		32'h00004554: begin
				q			<=			16'h2423;
		end
		32'h00004556: begin
				q			<=			16'h0CF1;
		end
		32'h00004558: begin
				q			<=			16'h0713;
		end
		32'h0000455A: begin
				q			<=			16'h0070;
		end
		32'h0000455C: begin
				q			<=			16'h8893;
		end
		32'h0000455E: begin
				q			<=			16'h0006;
		end
		32'h00004560: begin
				q			<=			16'h42E3;
		end
		32'h00004562: begin
				q			<=			16'hB4F7;
		end
		32'h00004564: begin
				q			<=			16'h7413;
		end
		32'h00004566: begin
				q			<=			16'h0044;
		end
		32'h00004568: begin
				q			<=			16'h1463;
		end
		32'h0000456A: begin
				q			<=			16'h7E04;
		end
		32'h0000456C: begin
				q			<=			16'h2D03;
		end
		32'h0000456E: begin
				q			<=			16'h01C1;
		end
		32'h00004570: begin
				q			<=			16'h2783;
		end
		32'h00004572: begin
				q			<=			16'h0201;
		end
		32'h00004574: begin
				q			<=			16'h5463;
		end
		32'h00004576: begin
				q			<=			16'h00FD;
		end
		32'h00004578: begin
				q			<=			16'h8D13;
		end
		32'h0000457A: begin
				q			<=			16'h0007;
		end
		32'h0000457C: begin
				q			<=			16'h2783;
		end
		32'h0000457E: begin
				q			<=			16'h0181;
		end
		32'h00004580: begin
				q			<=			16'h87B3;
		end
		32'h00004582: begin
				q			<=			16'h01A7;
		end
		32'h00004584: begin
				q			<=			16'h2C23;
		end
		32'h00004586: begin
				q			<=			16'h00F1;
		end
		32'h00004588: begin
				q			<=			16'h2783;
		end
		32'h0000458A: begin
				q			<=			16'h0CC1;
		end
		32'h0000458C: begin
				q			<=			16'h8C63;
		end
		32'h0000458E: begin
				q			<=			16'h0007;
		end
		32'h00004590: begin
				q			<=			16'h0613;
		end
		32'h00004592: begin
				q			<=			16'h0C41;
		end
		32'h00004594: begin
				q			<=			16'h8593;
		end
		32'h00004596: begin
				q			<=			16'h0009;
		end
		32'h00004598: begin
				q			<=			16'h0513;
		end
		32'h0000459A: begin
				q			<=			16'h0009;
		end
		32'h0000459C: begin
				q			<=			16'h40EF;
		end
		32'h0000459E: begin
				q			<=			16'h5C00;
		end
		32'h000045A0: begin
				q			<=			16'h18E3;
		end
		32'h000045A2: begin
				q			<=			16'h0005;
		end
		32'h000045A4: begin
				q			<=			16'h2783;
		end
		32'h000045A6: begin
				q			<=			16'h0041;
		end
		32'h000045A8: begin
				q			<=			16'h2423;
		end
		32'h000045AA: begin
				q			<=			16'h0C01;
		end
		32'h000045AC: begin
				q			<=			16'h9EE3;
		end
		32'h000045AE: begin
				q			<=			16'h0407;
		end
		32'h000045B0: begin
				q			<=			16'h0893;
		end
		32'h000045B2: begin
				q			<=			16'h0EC1;
		end
		32'h000045B4: begin
				q			<=			16'hF06F;
		end
		32'h000045B6: begin
				q			<=			16'hF14F;
		end
		32'h000045B8: begin
				q			<=			16'h0713;
		end
		32'h000045BA: begin
				q			<=			16'h0107;
		end
		32'h000045BC: begin
				q			<=			16'hA223;
		end
		32'h000045BE: begin
				q			<=			16'h0178;
		end
		32'h000045C0: begin
				q			<=			16'h2623;
		end
		32'h000045C2: begin
				q			<=			16'h0CE1;
		end
		32'h000045C4: begin
				q			<=			16'h2423;
		end
		32'h000045C6: begin
				q			<=			16'h0CF1;
		end
		32'h000045C8: begin
				q			<=			16'h5E63;
		end
		32'h000045CA: begin
				q			<=			16'h00FC;
		end
		32'h000045CC: begin
				q			<=			16'h0613;
		end
		32'h000045CE: begin
				q			<=			16'h0C41;
		end
		32'h000045D0: begin
				q			<=			16'h8593;
		end
		32'h000045D2: begin
				q			<=			16'h0009;
		end
		32'h000045D4: begin
				q			<=			16'h0513;
		end
		32'h000045D6: begin
				q			<=			16'h0009;
		end
		32'h000045D8: begin
				q			<=			16'h40EF;
		end
		32'h000045DA: begin
				q			<=			16'h5840;
		end
		32'h000045DC: begin
				q			<=			16'h1A63;
		end
		32'h000045DE: begin
				q			<=			16'h7C05;
		end
		32'h000045E0: begin
				q			<=			16'h0693;
		end
		32'h000045E2: begin
				q			<=			16'h0EC1;
		end
		32'h000045E4: begin
				q			<=			16'h8493;
		end
		32'h000045E6: begin
				q			<=			16'hFF04;
		end
		32'h000045E8: begin
				q			<=			16'h8893;
		end
		32'h000045EA: begin
				q			<=			16'h0006;
		end
		32'h000045EC: begin
				q			<=			16'hF06F;
		end
		32'h000045EE: begin
				q			<=			16'hF45F;
		end
		32'h000045F0: begin
				q			<=			16'h2703;
		end
		32'h000045F2: begin
				q			<=			16'h0AC1;
		end
		32'h000045F4: begin
				q			<=			16'h4663;
		end
		32'h000045F6: begin
				q			<=			16'h16E0;
		end
		32'h000045F8: begin
				q			<=			16'hB797;
		end
		32'h000045FA: begin
				q			<=			16'h0000;
		end
		32'h000045FC: begin
				q			<=			16'h8793;
		end
		32'h000045FE: begin
				q			<=			16'h7B47;
		end
		32'h00004600: begin
				q			<=			16'hA023;
		end
		32'h00004602: begin
				q			<=			16'h00F8;
		end
		32'h00004604: begin
				q			<=			16'h0793;
		end
		32'h00004606: begin
				q			<=			16'h0010;
		end
		32'h00004608: begin
				q			<=			16'hA223;
		end
		32'h0000460A: begin
				q			<=			16'h00F8;
		end
		32'h0000460C: begin
				q			<=			16'h2783;
		end
		32'h0000460E: begin
				q			<=			16'h0C81;
		end
		32'h00004610: begin
				q			<=			16'h8D93;
		end
		32'h00004612: begin
				q			<=			16'h001D;
		end
		32'h00004614: begin
				q			<=			16'h2623;
		end
		32'h00004616: begin
				q			<=			16'h0DB1;
		end
		32'h00004618: begin
				q			<=			16'h8793;
		end
		32'h0000461A: begin
				q			<=			16'h0017;
		end
		32'h0000461C: begin
				q			<=			16'h2423;
		end
		32'h0000461E: begin
				q			<=			16'h0CF1;
		end
		32'h00004620: begin
				q			<=			16'h0713;
		end
		32'h00004622: begin
				q			<=			16'h0070;
		end
		32'h00004624: begin
				q			<=			16'h8893;
		end
		32'h00004626: begin
				q			<=			16'h0088;
		end
		32'h00004628: begin
				q			<=			16'h5E63;
		end
		32'h0000462A: begin
				q			<=			16'h00F7;
		end
		32'h0000462C: begin
				q			<=			16'h0613;
		end
		32'h0000462E: begin
				q			<=			16'h0C41;
		end
		32'h00004630: begin
				q			<=			16'h8593;
		end
		32'h00004632: begin
				q			<=			16'h0009;
		end
		32'h00004634: begin
				q			<=			16'h0513;
		end
		32'h00004636: begin
				q			<=			16'h0009;
		end
		32'h00004638: begin
				q			<=			16'h40EF;
		end
		32'h0000463A: begin
				q			<=			16'h5240;
		end
		32'h0000463C: begin
				q			<=			16'h1A63;
		end
		32'h0000463E: begin
				q			<=			16'h7605;
		end
		32'h00004640: begin
				q			<=			16'h0893;
		end
		32'h00004642: begin
				q			<=			16'h0EC1;
		end
		32'h00004644: begin
				q			<=			16'h2783;
		end
		32'h00004646: begin
				q			<=			16'h0AC1;
		end
		32'h00004648: begin
				q			<=			16'h9863;
		end
		32'h0000464A: begin
				q			<=			16'h0007;
		end
		32'h0000464C: begin
				q			<=			16'h1663;
		end
		32'h0000464E: begin
				q			<=			16'h000A;
		end
		32'h00004650: begin
				q			<=			16'h7793;
		end
		32'h00004652: begin
				q			<=			16'h0014;
		end
		32'h00004654: begin
				q			<=			16'h88E3;
		end
		32'h00004656: begin
				q			<=			16'hF007;
		end
		32'h00004658: begin
				q			<=			16'h2783;
		end
		32'h0000465A: begin
				q			<=			16'h0281;
		end
		32'h0000465C: begin
				q			<=			16'h2703;
		end
		32'h0000465E: begin
				q			<=			16'h0141;
		end
		32'h00004660: begin
				q			<=			16'h8893;
		end
		32'h00004662: begin
				q			<=			16'h0088;
		end
		32'h00004664: begin
				q			<=			16'hAC23;
		end
		32'h00004666: begin
				q			<=			16'hFEF8;
		end
		32'h00004668: begin
				q			<=			16'h2783;
		end
		32'h0000466A: begin
				q			<=			16'h0141;
		end
		32'h0000466C: begin
				q			<=			16'hAE23;
		end
		32'h0000466E: begin
				q			<=			16'hFEF8;
		end
		32'h00004670: begin
				q			<=			16'h2783;
		end
		32'h00004672: begin
				q			<=			16'h0CC1;
		end
		32'h00004674: begin
				q			<=			16'h87B3;
		end
		32'h00004676: begin
				q			<=			16'h00E7;
		end
		32'h00004678: begin
				q			<=			16'h2623;
		end
		32'h0000467A: begin
				q			<=			16'h0CF1;
		end
		32'h0000467C: begin
				q			<=			16'h2783;
		end
		32'h0000467E: begin
				q			<=			16'h0C81;
		end
		32'h00004680: begin
				q			<=			16'h0713;
		end
		32'h00004682: begin
				q			<=			16'h0070;
		end
		32'h00004684: begin
				q			<=			16'h8793;
		end
		32'h00004686: begin
				q			<=			16'h0017;
		end
		32'h00004688: begin
				q			<=			16'h2423;
		end
		32'h0000468A: begin
				q			<=			16'h0CF1;
		end
		32'h0000468C: begin
				q			<=			16'h5E63;
		end
		32'h0000468E: begin
				q			<=			16'h00F7;
		end
		32'h00004690: begin
				q			<=			16'h0613;
		end
		32'h00004692: begin
				q			<=			16'h0C41;
		end
		32'h00004694: begin
				q			<=			16'h8593;
		end
		32'h00004696: begin
				q			<=			16'h0009;
		end
		32'h00004698: begin
				q			<=			16'h0513;
		end
		32'h0000469A: begin
				q			<=			16'h0009;
		end
		32'h0000469C: begin
				q			<=			16'h40EF;
		end
		32'h0000469E: begin
				q			<=			16'h4C00;
		end
		32'h000046A0: begin
				q			<=			16'h1863;
		end
		32'h000046A2: begin
				q			<=			16'h7005;
		end
		32'h000046A4: begin
				q			<=			16'h0893;
		end
		32'h000046A6: begin
				q			<=			16'h0EC1;
		end
		32'h000046A8: begin
				q			<=			16'h2A83;
		end
		32'h000046AA: begin
				q			<=			16'h0AC1;
		end
		32'h000046AC: begin
				q			<=			16'hD263;
		end
		32'h000046AE: begin
				q			<=			16'h060A;
		end
		32'h000046B0: begin
				q			<=			16'h0AB3;
		end
		32'h000046B2: begin
				q			<=			16'h4150;
		end
		32'h000046B4: begin
				q			<=			16'h8713;
		end
		32'h000046B6: begin
				q			<=			16'h0008;
		end
		32'h000046B8: begin
				q			<=			16'h0C13;
		end
		32'h000046BA: begin
				q			<=			16'h0100;
		end
		32'h000046BC: begin
				q			<=			16'hBB97;
		end
		32'h000046BE: begin
				q			<=			16'h0000;
		end
		32'h000046C0: begin
				q			<=			16'h8B93;
		end
		32'h000046C2: begin
				q			<=			16'hBE0B;
		end
		32'h000046C4: begin
				q			<=			16'h0D13;
		end
		32'h000046C6: begin
				q			<=			16'h0070;
		end
		32'h000046C8: begin
				q			<=			16'h2783;
		end
		32'h000046CA: begin
				q			<=			16'h0C81;
		end
		32'h000046CC: begin
				q			<=			16'h2023;
		end
		32'h000046CE: begin
				q			<=			16'h0177;
		end
		32'h000046D0: begin
				q			<=			16'h2683;
		end
		32'h000046D2: begin
				q			<=			16'h0CC1;
		end
		32'h000046D4: begin
				q			<=			16'h8793;
		end
		32'h000046D6: begin
				q			<=			16'h0017;
		end
		32'h000046D8: begin
				q			<=			16'h8893;
		end
		32'h000046DA: begin
				q			<=			16'h0088;
		end
		32'h000046DC: begin
				q			<=			16'h4663;
		end
		32'h000046DE: begin
				q			<=			16'h055C;
		end
		32'h000046E0: begin
				q			<=			16'h2223;
		end
		32'h000046E2: begin
				q			<=			16'h0157;
		end
		32'h000046E4: begin
				q			<=			16'h8AB3;
		end
		32'h000046E6: begin
				q			<=			16'h00DA;
		end
		32'h000046E8: begin
				q			<=			16'h2623;
		end
		32'h000046EA: begin
				q			<=			16'h0D51;
		end
		32'h000046EC: begin
				q			<=			16'h2423;
		end
		32'h000046EE: begin
				q			<=			16'h0CF1;
		end
		32'h000046F0: begin
				q			<=			16'h0713;
		end
		32'h000046F2: begin
				q			<=			16'h0070;
		end
		32'h000046F4: begin
				q			<=			16'h5E63;
		end
		32'h000046F6: begin
				q			<=			16'h00F7;
		end
		32'h000046F8: begin
				q			<=			16'h0613;
		end
		32'h000046FA: begin
				q			<=			16'h0C41;
		end
		32'h000046FC: begin
				q			<=			16'h8593;
		end
		32'h000046FE: begin
				q			<=			16'h0009;
		end
		32'h00004700: begin
				q			<=			16'h0513;
		end
		32'h00004702: begin
				q			<=			16'h0009;
		end
		32'h00004704: begin
				q			<=			16'h40EF;
		end
		32'h00004706: begin
				q			<=			16'h4580;
		end
		32'h00004708: begin
				q			<=			16'h1463;
		end
		32'h0000470A: begin
				q			<=			16'h6A05;
		end
		32'h0000470C: begin
				q			<=			16'h0893;
		end
		32'h0000470E: begin
				q			<=			16'h0EC1;
		end
		32'h00004710: begin
				q			<=			16'h2783;
		end
		32'h00004712: begin
				q			<=			16'h0CC1;
		end
		32'h00004714: begin
				q			<=			16'hA023;
		end
		32'h00004716: begin
				q			<=			16'h0098;
		end
		32'h00004718: begin
				q			<=			16'hA223;
		end
		32'h0000471A: begin
				q			<=			16'h0148;
		end
		32'h0000471C: begin
				q			<=			16'h87B3;
		end
		32'h0000471E: begin
				q			<=			16'h0147;
		end
		32'h00004720: begin
				q			<=			16'h2623;
		end
		32'h00004722: begin
				q			<=			16'h0CF1;
		end
		32'h00004724: begin
				q			<=			16'hF06F;
		end
		32'h00004726: begin
				q			<=			16'h969F;
		end
		32'h00004728: begin
				q			<=			16'h8693;
		end
		32'h0000472A: begin
				q			<=			16'h0106;
		end
		32'h0000472C: begin
				q			<=			16'h2223;
		end
		32'h0000472E: begin
				q			<=			16'h0187;
		end
		32'h00004730: begin
				q			<=			16'h2623;
		end
		32'h00004732: begin
				q			<=			16'h0CD1;
		end
		32'h00004734: begin
				q			<=			16'h2423;
		end
		32'h00004736: begin
				q			<=			16'h0CF1;
		end
		32'h00004738: begin
				q			<=			16'h5E63;
		end
		32'h0000473A: begin
				q			<=			16'h00FD;
		end
		32'h0000473C: begin
				q			<=			16'h0613;
		end
		32'h0000473E: begin
				q			<=			16'h0C41;
		end
		32'h00004740: begin
				q			<=			16'h8593;
		end
		32'h00004742: begin
				q			<=			16'h0009;
		end
		32'h00004744: begin
				q			<=			16'h0513;
		end
		32'h00004746: begin
				q			<=			16'h0009;
		end
		32'h00004748: begin
				q			<=			16'h40EF;
		end
		32'h0000474A: begin
				q			<=			16'h4140;
		end
		32'h0000474C: begin
				q			<=			16'h1263;
		end
		32'h0000474E: begin
				q			<=			16'h6605;
		end
		32'h00004750: begin
				q			<=			16'h0893;
		end
		32'h00004752: begin
				q			<=			16'h0EC1;
		end
		32'h00004754: begin
				q			<=			16'h8A93;
		end
		32'h00004756: begin
				q			<=			16'hFF0A;
		end
		32'h00004758: begin
				q			<=			16'h8713;
		end
		32'h0000475A: begin
				q			<=			16'h0008;
		end
		32'h0000475C: begin
				q			<=			16'hF06F;
		end
		32'h0000475E: begin
				q			<=			16'hF6DF;
		end
		32'h00004760: begin
				q			<=			16'h8A93;
		end
		32'h00004762: begin
				q			<=			16'h000C;
		end
		32'h00004764: begin
				q			<=			16'h5463;
		end
		32'h00004766: begin
				q			<=			16'h019A;
		end
		32'h00004768: begin
				q			<=			16'h0A93;
		end
		32'h0000476A: begin
				q			<=			16'h000A;
		end
		32'h0000476C: begin
				q			<=			16'h5263;
		end
		32'h0000476E: begin
				q			<=			16'h0550;
		end
		32'h00004770: begin
				q			<=			16'h2703;
		end
		32'h00004772: begin
				q			<=			16'h0C81;
		end
		32'h00004774: begin
				q			<=			16'h8DB3;
		end
		32'h00004776: begin
				q			<=			16'h01BA;
		end
		32'h00004778: begin
				q			<=			16'hA023;
		end
		32'h0000477A: begin
				q			<=			16'h0098;
		end
		32'h0000477C: begin
				q			<=			16'h0713;
		end
		32'h0000477E: begin
				q			<=			16'h0017;
		end
		32'h00004780: begin
				q			<=			16'hA223;
		end
		32'h00004782: begin
				q			<=			16'h0158;
		end
		32'h00004784: begin
				q			<=			16'h2623;
		end
		32'h00004786: begin
				q			<=			16'h0DB1;
		end
		32'h00004788: begin
				q			<=			16'h2423;
		end
		32'h0000478A: begin
				q			<=			16'h0CE1;
		end
		32'h0000478C: begin
				q			<=			16'h0693;
		end
		32'h0000478E: begin
				q			<=			16'h0070;
		end
		32'h00004790: begin
				q			<=			16'h8893;
		end
		32'h00004792: begin
				q			<=			16'h0088;
		end
		32'h00004794: begin
				q			<=			16'hDE63;
		end
		32'h00004796: begin
				q			<=			16'h00E6;
		end
		32'h00004798: begin
				q			<=			16'h0613;
		end
		32'h0000479A: begin
				q			<=			16'h0C41;
		end
		32'h0000479C: begin
				q			<=			16'h8593;
		end
		32'h0000479E: begin
				q			<=			16'h0009;
		end
		32'h000047A0: begin
				q			<=			16'h0513;
		end
		32'h000047A2: begin
				q			<=			16'h0009;
		end
		32'h000047A4: begin
				q			<=			16'h40EF;
		end
		32'h000047A6: begin
				q			<=			16'h3B80;
		end
		32'h000047A8: begin
				q			<=			16'h1463;
		end
		32'h000047AA: begin
				q			<=			16'h6005;
		end
		32'h000047AC: begin
				q			<=			16'h0893;
		end
		32'h000047AE: begin
				q			<=			16'h0EC1;
		end
		32'h000047B0: begin
				q			<=			16'hD463;
		end
		32'h000047B2: begin
				q			<=			16'h000A;
		end
		32'h000047B4: begin
				q			<=			16'h0A93;
		end
		32'h000047B6: begin
				q			<=			16'h0000;
		end
		32'h000047B8: begin
				q			<=			16'h8AB3;
		end
		32'h000047BA: begin
				q			<=			16'h415C;
		end
		32'h000047BC: begin
				q			<=			16'h5063;
		end
		32'h000047BE: begin
				q			<=			16'h0750;
		end
		32'h000047C0: begin
				q			<=			16'h0D93;
		end
		32'h000047C2: begin
				q			<=			16'h0100;
		end
		32'h000047C4: begin
				q			<=			16'hBD17;
		end
		32'h000047C6: begin
				q			<=			16'h0000;
		end
		32'h000047C8: begin
				q			<=			16'h0D13;
		end
		32'h000047CA: begin
				q			<=			16'hAD8D;
		end
		32'h000047CC: begin
				q			<=			16'h0B13;
		end
		32'h000047CE: begin
				q			<=			16'h0070;
		end
		32'h000047D0: begin
				q			<=			16'h2703;
		end
		32'h000047D2: begin
				q			<=			16'h0C81;
		end
		32'h000047D4: begin
				q			<=			16'hA023;
		end
		32'h000047D6: begin
				q			<=			16'h01A8;
		end
		32'h000047D8: begin
				q			<=			16'h2683;
		end
		32'h000047DA: begin
				q			<=			16'h0CC1;
		end
		32'h000047DC: begin
				q			<=			16'h0713;
		end
		32'h000047DE: begin
				q			<=			16'h0017;
		end
		32'h000047E0: begin
				q			<=			16'h8613;
		end
		32'h000047E2: begin
				q			<=			16'h0088;
		end
		32'h000047E4: begin
				q			<=			16'hC263;
		end
		32'h000047E6: begin
				q			<=			16'h1B5D;
		end
		32'h000047E8: begin
				q			<=			16'hA223;
		end
		32'h000047EA: begin
				q			<=			16'h0158;
		end
		32'h000047EC: begin
				q			<=			16'h8AB3;
		end
		32'h000047EE: begin
				q			<=			16'h00DA;
		end
		32'h000047F0: begin
				q			<=			16'h2623;
		end
		32'h000047F2: begin
				q			<=			16'h0D51;
		end
		32'h000047F4: begin
				q			<=			16'h2423;
		end
		32'h000047F6: begin
				q			<=			16'h0CE1;
		end
		32'h000047F8: begin
				q			<=			16'h0693;
		end
		32'h000047FA: begin
				q			<=			16'h0070;
		end
		32'h000047FC: begin
				q			<=			16'h0893;
		end
		32'h000047FE: begin
				q			<=			16'h0006;
		end
		32'h00004800: begin
				q			<=			16'hDE63;
		end
		32'h00004802: begin
				q			<=			16'h00E6;
		end
		32'h00004804: begin
				q			<=			16'h0613;
		end
		32'h00004806: begin
				q			<=			16'h0C41;
		end
		32'h00004808: begin
				q			<=			16'h8593;
		end
		32'h0000480A: begin
				q			<=			16'h0009;
		end
		32'h0000480C: begin
				q			<=			16'h0513;
		end
		32'h0000480E: begin
				q			<=			16'h0009;
		end
		32'h00004810: begin
				q			<=			16'h40EF;
		end
		32'h00004812: begin
				q			<=			16'h34C0;
		end
		32'h00004814: begin
				q			<=			16'h1E63;
		end
		32'h00004816: begin
				q			<=			16'h5805;
		end
		32'h00004818: begin
				q			<=			16'h0893;
		end
		32'h0000481A: begin
				q			<=			16'h0EC1;
		end
		32'h0000481C: begin
				q			<=			16'h7793;
		end
		32'h0000481E: begin
				q			<=			16'h4004;
		end
		32'h00004820: begin
				q			<=			16'h8AB3;
		end
		32'h00004822: begin
				q			<=			16'h0194;
		end
		32'h00004824: begin
				q			<=			16'h8463;
		end
		32'h00004826: begin
				q			<=			16'h0207;
		end
		32'h00004828: begin
				q			<=			16'h0D13;
		end
		32'h0000482A: begin
				q			<=			16'h0070;
		end
		32'h0000482C: begin
				q			<=			16'h8B33;
		end
		32'h0000482E: begin
				q			<=			16'h0144;
		end
		32'h00004830: begin
				q			<=			16'hBD97;
		end
		32'h00004832: begin
				q			<=			16'h0000;
		end
		32'h00004834: begin
				q			<=			16'h8D93;
		end
		32'h00004836: begin
				q			<=			16'hA6CD;
		end
		32'h00004838: begin
				q			<=			16'h9463;
		end
		32'h0000483A: begin
				q			<=			16'h180B;
		end
		32'h0000483C: begin
				q			<=			16'h1463;
		end
		32'h0000483E: begin
				q			<=			16'h180C;
		end
		32'h00004840: begin
				q			<=			16'h87B3;
		end
		32'h00004842: begin
				q			<=			16'h0144;
		end
		32'h00004844: begin
				q			<=			16'hF463;
		end
		32'h00004846: begin
				q			<=			16'h0157;
		end
		32'h00004848: begin
				q			<=			16'h8A93;
		end
		32'h0000484A: begin
				q			<=			16'h0007;
		end
		32'h0000484C: begin
				q			<=			16'h2783;
		end
		32'h0000484E: begin
				q			<=			16'h0AC1;
		end
		32'h00004850: begin
				q			<=			16'hC663;
		end
		32'h00004852: begin
				q			<=			16'h0147;
		end
		32'h00004854: begin
				q			<=			16'h7793;
		end
		32'h00004856: begin
				q			<=			16'h0014;
		end
		32'h00004858: begin
				q			<=			16'h8A63;
		end
		32'h0000485A: begin
				q			<=			16'h0407;
		end
		32'h0000485C: begin
				q			<=			16'h2783;
		end
		32'h0000485E: begin
				q			<=			16'h0281;
		end
		32'h00004860: begin
				q			<=			16'h2703;
		end
		32'h00004862: begin
				q			<=			16'h0141;
		end
		32'h00004864: begin
				q			<=			16'h8893;
		end
		32'h00004866: begin
				q			<=			16'h0088;
		end
		32'h00004868: begin
				q			<=			16'hAC23;
		end
		32'h0000486A: begin
				q			<=			16'hFEF8;
		end
		32'h0000486C: begin
				q			<=			16'h2783;
		end
		32'h0000486E: begin
				q			<=			16'h0141;
		end
		32'h00004870: begin
				q			<=			16'hAE23;
		end
		32'h00004872: begin
				q			<=			16'hFEF8;
		end
		32'h00004874: begin
				q			<=			16'h2783;
		end
		32'h00004876: begin
				q			<=			16'h0CC1;
		end
		32'h00004878: begin
				q			<=			16'h87B3;
		end
		32'h0000487A: begin
				q			<=			16'h00E7;
		end
		32'h0000487C: begin
				q			<=			16'h2623;
		end
		32'h0000487E: begin
				q			<=			16'h0CF1;
		end
		32'h00004880: begin
				q			<=			16'h2783;
		end
		32'h00004882: begin
				q			<=			16'h0C81;
		end
		32'h00004884: begin
				q			<=			16'h0713;
		end
		32'h00004886: begin
				q			<=			16'h0070;
		end
		32'h00004888: begin
				q			<=			16'h8793;
		end
		32'h0000488A: begin
				q			<=			16'h0017;
		end
		32'h0000488C: begin
				q			<=			16'h2423;
		end
		32'h0000488E: begin
				q			<=			16'h0CF1;
		end
		32'h00004890: begin
				q			<=			16'h5E63;
		end
		32'h00004892: begin
				q			<=			16'h00F7;
		end
		32'h00004894: begin
				q			<=			16'h0613;
		end
		32'h00004896: begin
				q			<=			16'h0C41;
		end
		32'h00004898: begin
				q			<=			16'h8593;
		end
		32'h0000489A: begin
				q			<=			16'h0009;
		end
		32'h0000489C: begin
				q			<=			16'h0513;
		end
		32'h0000489E: begin
				q			<=			16'h0009;
		end
		32'h000048A0: begin
				q			<=			16'h40EF;
		end
		32'h000048A2: begin
				q			<=			16'h2BC0;
		end
		32'h000048A4: begin
				q			<=			16'h1663;
		end
		32'h000048A6: begin
				q			<=			16'h5005;
		end
		32'h000048A8: begin
				q			<=			16'h0893;
		end
		32'h000048AA: begin
				q			<=			16'h0EC1;
		end
		32'h000048AC: begin
				q			<=			16'h84B3;
		end
		32'h000048AE: begin
				q			<=			16'h0144;
		end
		32'h000048B0: begin
				q			<=			16'h87B3;
		end
		32'h000048B2: begin
				q			<=			16'h4154;
		end
		32'h000048B4: begin
				q			<=			16'h2483;
		end
		32'h000048B6: begin
				q			<=			16'h0AC1;
		end
		32'h000048B8: begin
				q			<=			16'h04B3;
		end
		32'h000048BA: begin
				q			<=			16'h409A;
		end
		32'h000048BC: begin
				q			<=			16'hD463;
		end
		32'h000048BE: begin
				q			<=			16'h0097;
		end
		32'h000048C0: begin
				q			<=			16'h8493;
		end
		32'h000048C2: begin
				q			<=			16'h0007;
		end
		32'h000048C4: begin
				q			<=			16'h5463;
		end
		32'h000048C6: begin
				q			<=			16'h0490;
		end
		32'h000048C8: begin
				q			<=			16'h2783;
		end
		32'h000048CA: begin
				q			<=			16'h0CC1;
		end
		32'h000048CC: begin
				q			<=			16'hA023;
		end
		32'h000048CE: begin
				q			<=			16'h0158;
		end
		32'h000048D0: begin
				q			<=			16'hA223;
		end
		32'h000048D2: begin
				q			<=			16'h0098;
		end
		32'h000048D4: begin
				q			<=			16'h87B3;
		end
		32'h000048D6: begin
				q			<=			16'h00F4;
		end
		32'h000048D8: begin
				q			<=			16'h2623;
		end
		32'h000048DA: begin
				q			<=			16'h0CF1;
		end
		32'h000048DC: begin
				q			<=			16'h2783;
		end
		32'h000048DE: begin
				q			<=			16'h0C81;
		end
		32'h000048E0: begin
				q			<=			16'h0713;
		end
		32'h000048E2: begin
				q			<=			16'h0070;
		end
		32'h000048E4: begin
				q			<=			16'h8893;
		end
		32'h000048E6: begin
				q			<=			16'h0088;
		end
		32'h000048E8: begin
				q			<=			16'h8793;
		end
		32'h000048EA: begin
				q			<=			16'h0017;
		end
		32'h000048EC: begin
				q			<=			16'h2423;
		end
		32'h000048EE: begin
				q			<=			16'h0CF1;
		end
		32'h000048F0: begin
				q			<=			16'h5E63;
		end
		32'h000048F2: begin
				q			<=			16'h00F7;
		end
		32'h000048F4: begin
				q			<=			16'h0613;
		end
		32'h000048F6: begin
				q			<=			16'h0C41;
		end
		32'h000048F8: begin
				q			<=			16'h8593;
		end
		32'h000048FA: begin
				q			<=			16'h0009;
		end
		32'h000048FC: begin
				q			<=			16'h0513;
		end
		32'h000048FE: begin
				q			<=			16'h0009;
		end
		32'h00004900: begin
				q			<=			16'h40EF;
		end
		32'h00004902: begin
				q			<=			16'h25C0;
		end
		32'h00004904: begin
				q			<=			16'h1663;
		end
		32'h00004906: begin
				q			<=			16'h4A05;
		end
		32'h00004908: begin
				q			<=			16'h0893;
		end
		32'h0000490A: begin
				q			<=			16'h0EC1;
		end
		32'h0000490C: begin
				q			<=			16'h8793;
		end
		32'h0000490E: begin
				q			<=			16'h0004;
		end
		32'h00004910: begin
				q			<=			16'hD463;
		end
		32'h00004912: begin
				q			<=			16'h0004;
		end
		32'h00004914: begin
				q			<=			16'h0793;
		end
		32'h00004916: begin
				q			<=			16'h0000;
		end
		32'h00004918: begin
				q			<=			16'h2483;
		end
		32'h0000491A: begin
				q			<=			16'h0AC1;
		end
		32'h0000491C: begin
				q			<=			16'h04B3;
		end
		32'h0000491E: begin
				q			<=			16'h409A;
		end
		32'h00004920: begin
				q			<=			16'h84B3;
		end
		32'h00004922: begin
				q			<=			16'h40F4;
		end
		32'h00004924: begin
				q			<=			16'h50E3;
		end
		32'h00004926: begin
				q			<=			16'hC490;
		end
		32'h00004928: begin
				q			<=			16'h0B93;
		end
		32'h0000492A: begin
				q			<=			16'h0100;
		end
		32'h0000492C: begin
				q			<=			16'hBA97;
		end
		32'h0000492E: begin
				q			<=			16'h0000;
		end
		32'h00004930: begin
				q			<=			16'h8A93;
		end
		32'h00004932: begin
				q			<=			16'h970A;
		end
		32'h00004934: begin
				q			<=			16'h0C13;
		end
		32'h00004936: begin
				q			<=			16'h0070;
		end
		32'h00004938: begin
				q			<=			16'h2783;
		end
		32'h0000493A: begin
				q			<=			16'h0C81;
		end
		32'h0000493C: begin
				q			<=			16'hA023;
		end
		32'h0000493E: begin
				q			<=			16'h0158;
		end
		32'h00004940: begin
				q			<=			16'h2703;
		end
		32'h00004942: begin
				q			<=			16'h0CC1;
		end
		32'h00004944: begin
				q			<=			16'h8793;
		end
		32'h00004946: begin
				q			<=			16'h0017;
		end
		32'h00004948: begin
				q			<=			16'h8693;
		end
		32'h0000494A: begin
				q			<=			16'h0088;
		end
		32'h0000494C: begin
				q			<=			16'hDEE3;
		end
		32'h0000494E: begin
				q			<=			16'hBE9B;
		end
		32'h00004950: begin
				q			<=			16'h0713;
		end
		32'h00004952: begin
				q			<=			16'h0107;
		end
		32'h00004954: begin
				q			<=			16'hA223;
		end
		32'h00004956: begin
				q			<=			16'h0178;
		end
		32'h00004958: begin
				q			<=			16'h2623;
		end
		32'h0000495A: begin
				q			<=			16'h0CE1;
		end
		32'h0000495C: begin
				q			<=			16'h2423;
		end
		32'h0000495E: begin
				q			<=			16'h0CF1;
		end
		32'h00004960: begin
				q			<=			16'h5E63;
		end
		32'h00004962: begin
				q			<=			16'h00FC;
		end
		32'h00004964: begin
				q			<=			16'h0613;
		end
		32'h00004966: begin
				q			<=			16'h0C41;
		end
		32'h00004968: begin
				q			<=			16'h8593;
		end
		32'h0000496A: begin
				q			<=			16'h0009;
		end
		32'h0000496C: begin
				q			<=			16'h0513;
		end
		32'h0000496E: begin
				q			<=			16'h0009;
		end
		32'h00004970: begin
				q			<=			16'h40EF;
		end
		32'h00004972: begin
				q			<=			16'h1EC0;
		end
		32'h00004974: begin
				q			<=			16'h1E63;
		end
		32'h00004976: begin
				q			<=			16'h4205;
		end
		32'h00004978: begin
				q			<=			16'h0693;
		end
		32'h0000497A: begin
				q			<=			16'h0EC1;
		end
		32'h0000497C: begin
				q			<=			16'h8493;
		end
		32'h0000497E: begin
				q			<=			16'hFF04;
		end
		32'h00004980: begin
				q			<=			16'h8893;
		end
		32'h00004982: begin
				q			<=			16'h0006;
		end
		32'h00004984: begin
				q			<=			16'hF06F;
		end
		32'h00004986: begin
				q			<=			16'hFB5F;
		end
		32'h00004988: begin
				q			<=			16'h8693;
		end
		32'h0000498A: begin
				q			<=			16'h0106;
		end
		32'h0000498C: begin
				q			<=			16'hA223;
		end
		32'h0000498E: begin
				q			<=			16'h01B8;
		end
		32'h00004990: begin
				q			<=			16'h2623;
		end
		32'h00004992: begin
				q			<=			16'h0CD1;
		end
		32'h00004994: begin
				q			<=			16'h2423;
		end
		32'h00004996: begin
				q			<=			16'h0CE1;
		end
		32'h00004998: begin
				q			<=			16'h5E63;
		end
		32'h0000499A: begin
				q			<=			16'h00EB;
		end
		32'h0000499C: begin
				q			<=			16'h0613;
		end
		32'h0000499E: begin
				q			<=			16'h0C41;
		end
		32'h000049A0: begin
				q			<=			16'h8593;
		end
		32'h000049A2: begin
				q			<=			16'h0009;
		end
		32'h000049A4: begin
				q			<=			16'h0513;
		end
		32'h000049A6: begin
				q			<=			16'h0009;
		end
		32'h000049A8: begin
				q			<=			16'h40EF;
		end
		32'h000049AA: begin
				q			<=			16'h1B40;
		end
		32'h000049AC: begin
				q			<=			16'h1263;
		end
		32'h000049AE: begin
				q			<=			16'h4005;
		end
		32'h000049B0: begin
				q			<=			16'h0613;
		end
		32'h000049B2: begin
				q			<=			16'h0EC1;
		end
		32'h000049B4: begin
				q			<=			16'h8A93;
		end
		32'h000049B6: begin
				q			<=			16'hFF0A;
		end
		32'h000049B8: begin
				q			<=			16'h0893;
		end
		32'h000049BA: begin
				q			<=			16'h0006;
		end
		32'h000049BC: begin
				q			<=			16'hF06F;
		end
		32'h000049BE: begin
				q			<=			16'hE15F;
		end
		32'h000049C0: begin
				q			<=			16'h0263;
		end
		32'h000049C2: begin
				q			<=			16'h0E0C;
		end
		32'h000049C4: begin
				q			<=			16'h0C13;
		end
		32'h000049C6: begin
				q			<=			16'hFFFC;
		end
		32'h000049C8: begin
				q			<=			16'h2783;
		end
		32'h000049CA: begin
				q			<=			16'h02C1;
		end
		32'h000049CC: begin
				q			<=			16'h2703;
		end
		32'h000049CE: begin
				q			<=			16'h0241;
		end
		32'h000049D0: begin
				q			<=			16'h8893;
		end
		32'h000049D2: begin
				q			<=			16'h0088;
		end
		32'h000049D4: begin
				q			<=			16'hAC23;
		end
		32'h000049D6: begin
				q			<=			16'hFEF8;
		end
		32'h000049D8: begin
				q			<=			16'h2783;
		end
		32'h000049DA: begin
				q			<=			16'h0241;
		end
		32'h000049DC: begin
				q			<=			16'hAE23;
		end
		32'h000049DE: begin
				q			<=			16'hFEF8;
		end
		32'h000049E0: begin
				q			<=			16'h2783;
		end
		32'h000049E2: begin
				q			<=			16'h0CC1;
		end
		32'h000049E4: begin
				q			<=			16'h87B3;
		end
		32'h000049E6: begin
				q			<=			16'h00E7;
		end
		32'h000049E8: begin
				q			<=			16'h2623;
		end
		32'h000049EA: begin
				q			<=			16'h0CF1;
		end
		32'h000049EC: begin
				q			<=			16'h2783;
		end
		32'h000049EE: begin
				q			<=			16'h0C81;
		end
		32'h000049F0: begin
				q			<=			16'h8793;
		end
		32'h000049F2: begin
				q			<=			16'h0017;
		end
		32'h000049F4: begin
				q			<=			16'h2423;
		end
		32'h000049F6: begin
				q			<=			16'h0CF1;
		end
		32'h000049F8: begin
				q			<=			16'h5E63;
		end
		32'h000049FA: begin
				q			<=			16'h00FD;
		end
		32'h000049FC: begin
				q			<=			16'h0613;
		end
		32'h000049FE: begin
				q			<=			16'h0C41;
		end
		32'h00004A00: begin
				q			<=			16'h8593;
		end
		32'h00004A02: begin
				q			<=			16'h0009;
		end
		32'h00004A04: begin
				q			<=			16'h0513;
		end
		32'h00004A06: begin
				q			<=			16'h0009;
		end
		32'h00004A08: begin
				q			<=			16'h40EF;
		end
		32'h00004A0A: begin
				q			<=			16'h1540;
		end
		32'h00004A0C: begin
				q			<=			16'h1263;
		end
		32'h00004A0E: begin
				q			<=			16'h3A05;
		end
		32'h00004A10: begin
				q			<=			16'h0893;
		end
		32'h00004A12: begin
				q			<=			16'h0EC1;
		end
		32'h00004A14: begin
				q			<=			16'h2783;
		end
		32'h00004A16: begin
				q			<=			16'h0081;
		end
		32'h00004A18: begin
				q			<=			16'h0733;
		end
		32'h00004A1A: begin
				q			<=			16'h415B;
		end
		32'h00004A1C: begin
				q			<=			16'hC783;
		end
		32'h00004A1E: begin
				q			<=			16'h0007;
		end
		32'h00004A20: begin
				q			<=			16'h5463;
		end
		32'h00004A22: begin
				q			<=			16'h00F7;
		end
		32'h00004A24: begin
				q			<=			16'h0793;
		end
		32'h00004A26: begin
				q			<=			16'h0007;
		end
		32'h00004A28: begin
				q			<=			16'h5663;
		end
		32'h00004A2A: begin
				q			<=			16'h04F0;
		end
		32'h00004A2C: begin
				q			<=			16'h2703;
		end
		32'h00004A2E: begin
				q			<=			16'h0CC1;
		end
		32'h00004A30: begin
				q			<=			16'hA023;
		end
		32'h00004A32: begin
				q			<=			16'h0158;
		end
		32'h00004A34: begin
				q			<=			16'hA223;
		end
		32'h00004A36: begin
				q			<=			16'h00F8;
		end
		32'h00004A38: begin
				q			<=			16'h8733;
		end
		32'h00004A3A: begin
				q			<=			16'h00E7;
		end
		32'h00004A3C: begin
				q			<=			16'h2623;
		end
		32'h00004A3E: begin
				q			<=			16'h0CE1;
		end
		32'h00004A40: begin
				q			<=			16'h2703;
		end
		32'h00004A42: begin
				q			<=			16'h0C81;
		end
		32'h00004A44: begin
				q			<=			16'h8893;
		end
		32'h00004A46: begin
				q			<=			16'h0088;
		end
		32'h00004A48: begin
				q			<=			16'h0713;
		end
		32'h00004A4A: begin
				q			<=			16'h0017;
		end
		32'h00004A4C: begin
				q			<=			16'h2423;
		end
		32'h00004A4E: begin
				q			<=			16'h0CE1;
		end
		32'h00004A50: begin
				q			<=			16'h5263;
		end
		32'h00004A52: begin
				q			<=			16'h02ED;
		end
		32'h00004A54: begin
				q			<=			16'h0613;
		end
		32'h00004A56: begin
				q			<=			16'h0C41;
		end
		32'h00004A58: begin
				q			<=			16'h8593;
		end
		32'h00004A5A: begin
				q			<=			16'h0009;
		end
		32'h00004A5C: begin
				q			<=			16'h0513;
		end
		32'h00004A5E: begin
				q			<=			16'h0009;
		end
		32'h00004A60: begin
				q			<=			16'h2C23;
		end
		32'h00004A62: begin
				q			<=			16'h02F1;
		end
		32'h00004A64: begin
				q			<=			16'h40EF;
		end
		32'h00004A66: begin
				q			<=			16'h0F80;
		end
		32'h00004A68: begin
				q			<=			16'h1463;
		end
		32'h00004A6A: begin
				q			<=			16'h3405;
		end
		32'h00004A6C: begin
				q			<=			16'h2783;
		end
		32'h00004A6E: begin
				q			<=			16'h0381;
		end
		32'h00004A70: begin
				q			<=			16'h0893;
		end
		32'h00004A72: begin
				q			<=			16'h0EC1;
		end
		32'h00004A74: begin
				q			<=			16'h8713;
		end
		32'h00004A76: begin
				q			<=			16'h0007;
		end
		32'h00004A78: begin
				q			<=			16'hD463;
		end
		32'h00004A7A: begin
				q			<=			16'h0007;
		end
		32'h00004A7C: begin
				q			<=			16'h0713;
		end
		32'h00004A7E: begin
				q			<=			16'h0000;
		end
		32'h00004A80: begin
				q			<=			16'h2783;
		end
		32'h00004A82: begin
				q			<=			16'h0081;
		end
		32'h00004A84: begin
				q			<=			16'h0813;
		end
		32'h00004A86: begin
				q			<=			16'h0100;
		end
		32'h00004A88: begin
				q			<=			16'hC783;
		end
		32'h00004A8A: begin
				q			<=			16'h0007;
		end
		32'h00004A8C: begin
				q			<=			16'h87B3;
		end
		32'h00004A8E: begin
				q			<=			16'h40E7;
		end
		32'h00004A90: begin
				q			<=			16'h4663;
		end
		32'h00004A92: begin
				q			<=			16'h06F0;
		end
		32'h00004A94: begin
				q			<=			16'h2783;
		end
		32'h00004A96: begin
				q			<=			16'h0081;
		end
		32'h00004A98: begin
				q			<=			16'hC783;
		end
		32'h00004A9A: begin
				q			<=			16'h0007;
		end
		32'h00004A9C: begin
				q			<=			16'h8AB3;
		end
		32'h00004A9E: begin
				q			<=			16'h00FA;
		end
		32'h00004AA0: begin
				q			<=			16'hF06F;
		end
		32'h00004AA2: begin
				q			<=			16'hD99F;
		end
		32'h00004AA4: begin
				q			<=			16'h2783;
		end
		32'h00004AA6: begin
				q			<=			16'h0081;
		end
		32'h00004AA8: begin
				q			<=			16'h8B93;
		end
		32'h00004AAA: begin
				q			<=			16'hFFFB;
		end
		32'h00004AAC: begin
				q			<=			16'h8793;
		end
		32'h00004AAE: begin
				q			<=			16'hFFF7;
		end
		32'h00004AB0: begin
				q			<=			16'h2423;
		end
		32'h00004AB2: begin
				q			<=			16'h00F1;
		end
		32'h00004AB4: begin
				q			<=			16'hF06F;
		end
		32'h00004AB6: begin
				q			<=			16'hF15F;
		end
		32'h00004AB8: begin
				q			<=			16'h8693;
		end
		32'h00004ABA: begin
				q			<=			16'h0106;
		end
		32'h00004ABC: begin
				q			<=			16'hA223;
		end
		32'h00004ABE: begin
				q			<=			16'h0108;
		end
		32'h00004AC0: begin
				q			<=			16'h2623;
		end
		32'h00004AC2: begin
				q			<=			16'h0CD1;
		end
		32'h00004AC4: begin
				q			<=			16'h2423;
		end
		32'h00004AC6: begin
				q			<=			16'h0CE1;
		end
		32'h00004AC8: begin
				q			<=			16'h5663;
		end
		32'h00004ACA: begin
				q			<=			16'h02ED;
		end
		32'h00004ACC: begin
				q			<=			16'h0613;
		end
		32'h00004ACE: begin
				q			<=			16'h0C41;
		end
		32'h00004AD0: begin
				q			<=			16'h8593;
		end
		32'h00004AD2: begin
				q			<=			16'h0009;
		end
		32'h00004AD4: begin
				q			<=			16'h0513;
		end
		32'h00004AD6: begin
				q			<=			16'h0009;
		end
		32'h00004AD8: begin
				q			<=			16'h2E23;
		end
		32'h00004ADA: begin
				q			<=			16'h0301;
		end
		32'h00004ADC: begin
				q			<=			16'h2C23;
		end
		32'h00004ADE: begin
				q			<=			16'h02F1;
		end
		32'h00004AE0: begin
				q			<=			16'h40EF;
		end
		32'h00004AE2: begin
				q			<=			16'h07C0;
		end
		32'h00004AE4: begin
				q			<=			16'h1663;
		end
		32'h00004AE6: begin
				q			<=			16'h2C05;
		end
		32'h00004AE8: begin
				q			<=			16'h2803;
		end
		32'h00004AEA: begin
				q			<=			16'h03C1;
		end
		32'h00004AEC: begin
				q			<=			16'h2783;
		end
		32'h00004AEE: begin
				q			<=			16'h0381;
		end
		32'h00004AF0: begin
				q			<=			16'h0613;
		end
		32'h00004AF2: begin
				q			<=			16'h0EC1;
		end
		32'h00004AF4: begin
				q			<=			16'h8793;
		end
		32'h00004AF6: begin
				q			<=			16'hFF07;
		end
		32'h00004AF8: begin
				q			<=			16'h0893;
		end
		32'h00004AFA: begin
				q			<=			16'h0006;
		end
		32'h00004AFC: begin
				q			<=			16'h2703;
		end
		32'h00004AFE: begin
				q			<=			16'h0C81;
		end
		32'h00004B00: begin
				q			<=			16'hA023;
		end
		32'h00004B02: begin
				q			<=			16'h01B8;
		end
		32'h00004B04: begin
				q			<=			16'h2683;
		end
		32'h00004B06: begin
				q			<=			16'h0CC1;
		end
		32'h00004B08: begin
				q			<=			16'h0713;
		end
		32'h00004B0A: begin
				q			<=			16'h0017;
		end
		32'h00004B0C: begin
				q			<=			16'h8613;
		end
		32'h00004B0E: begin
				q			<=			16'h0088;
		end
		32'h00004B10: begin
				q			<=			16'h44E3;
		end
		32'h00004B12: begin
				q			<=			16'hFAF8;
		end
		32'h00004B14: begin
				q			<=			16'hA223;
		end
		32'h00004B16: begin
				q			<=			16'h00F8;
		end
		32'h00004B18: begin
				q			<=			16'h87B3;
		end
		32'h00004B1A: begin
				q			<=			16'h00D7;
		end
		32'h00004B1C: begin
				q			<=			16'h2623;
		end
		32'h00004B1E: begin
				q			<=			16'h0CF1;
		end
		32'h00004B20: begin
				q			<=			16'h2423;
		end
		32'h00004B22: begin
				q			<=			16'h0CE1;
		end
		32'h00004B24: begin
				q			<=			16'h0893;
		end
		32'h00004B26: begin
				q			<=			16'h0006;
		end
		32'h00004B28: begin
				q			<=			16'h56E3;
		end
		32'h00004B2A: begin
				q			<=			16'hF6ED;
		end
		32'h00004B2C: begin
				q			<=			16'h0613;
		end
		32'h00004B2E: begin
				q			<=			16'h0C41;
		end
		32'h00004B30: begin
				q			<=			16'h8593;
		end
		32'h00004B32: begin
				q			<=			16'h0009;
		end
		32'h00004B34: begin
				q			<=			16'h0513;
		end
		32'h00004B36: begin
				q			<=			16'h0009;
		end
		32'h00004B38: begin
				q			<=			16'h40EF;
		end
		32'h00004B3A: begin
				q			<=			16'h0240;
		end
		32'h00004B3C: begin
				q			<=			16'h1A63;
		end
		32'h00004B3E: begin
				q			<=			16'h2605;
		end
		32'h00004B40: begin
				q			<=			16'h0893;
		end
		32'h00004B42: begin
				q			<=			16'h0EC1;
		end
		32'h00004B44: begin
				q			<=			16'hF06F;
		end
		32'h00004B46: begin
				q			<=			16'hF51F;
		end
		32'h00004B48: begin
				q			<=			16'h2783;
		end
		32'h00004B4A: begin
				q			<=			16'h0C81;
		end
		32'h00004B4C: begin
				q			<=			16'h0713;
		end
		32'h00004B4E: begin
				q			<=			16'h0010;
		end
		32'h00004B50: begin
				q			<=			16'hA023;
		end
		32'h00004B52: begin
				q			<=			16'h0098;
		end
		32'h00004B54: begin
				q			<=			16'h8D93;
		end
		32'h00004B56: begin
				q			<=			16'h001D;
		end
		32'h00004B58: begin
				q			<=			16'h8793;
		end
		32'h00004B5A: begin
				q			<=			16'h0017;
		end
		32'h00004B5C: begin
				q			<=			16'h8B93;
		end
		32'h00004B5E: begin
				q			<=			16'h0088;
		end
		32'h00004B60: begin
				q			<=			16'h4663;
		end
		32'h00004B62: begin
				q			<=			16'h0147;
		end
		32'h00004B64: begin
				q			<=			16'h7693;
		end
		32'h00004B66: begin
				q			<=			16'h0014;
		end
		32'h00004B68: begin
				q			<=			16'h8863;
		end
		32'h00004B6A: begin
				q			<=			16'h1C06;
		end
		32'h00004B6C: begin
				q			<=			16'h0713;
		end
		32'h00004B6E: begin
				q			<=			16'h0010;
		end
		32'h00004B70: begin
				q			<=			16'hA223;
		end
		32'h00004B72: begin
				q			<=			16'h00E8;
		end
		32'h00004B74: begin
				q			<=			16'h2623;
		end
		32'h00004B76: begin
				q			<=			16'h0DB1;
		end
		32'h00004B78: begin
				q			<=			16'h2423;
		end
		32'h00004B7A: begin
				q			<=			16'h0CF1;
		end
		32'h00004B7C: begin
				q			<=			16'h0713;
		end
		32'h00004B7E: begin
				q			<=			16'h0070;
		end
		32'h00004B80: begin
				q			<=			16'h5E63;
		end
		32'h00004B82: begin
				q			<=			16'h00F7;
		end
		32'h00004B84: begin
				q			<=			16'h0613;
		end
		32'h00004B86: begin
				q			<=			16'h0C41;
		end
		32'h00004B88: begin
				q			<=			16'h8593;
		end
		32'h00004B8A: begin
				q			<=			16'h0009;
		end
		32'h00004B8C: begin
				q			<=			16'h0513;
		end
		32'h00004B8E: begin
				q			<=			16'h0009;
		end
		32'h00004B90: begin
				q			<=			16'h30EF;
		end
		32'h00004B92: begin
				q			<=			16'h7CD0;
		end
		32'h00004B94: begin
				q			<=			16'h1E63;
		end
		32'h00004B96: begin
				q			<=			16'h2005;
		end
		32'h00004B98: begin
				q			<=			16'h0B93;
		end
		32'h00004B9A: begin
				q			<=			16'h0EC1;
		end
		32'h00004B9C: begin
				q			<=			16'h2783;
		end
		32'h00004B9E: begin
				q			<=			16'h0281;
		end
		32'h00004BA0: begin
				q			<=			16'h2703;
		end
		32'h00004BA2: begin
				q			<=			16'h0141;
		end
		32'h00004BA4: begin
				q			<=			16'h8B93;
		end
		32'h00004BA6: begin
				q			<=			16'h008B;
		end
		32'h00004BA8: begin
				q			<=			16'hAC23;
		end
		32'h00004BAA: begin
				q			<=			16'hFEFB;
		end
		32'h00004BAC: begin
				q			<=			16'h2783;
		end
		32'h00004BAE: begin
				q			<=			16'h0141;
		end
		32'h00004BB0: begin
				q			<=			16'hAE23;
		end
		32'h00004BB2: begin
				q			<=			16'hFEFB;
		end
		32'h00004BB4: begin
				q			<=			16'h2783;
		end
		32'h00004BB6: begin
				q			<=			16'h0CC1;
		end
		32'h00004BB8: begin
				q			<=			16'h87B3;
		end
		32'h00004BBA: begin
				q			<=			16'h00E7;
		end
		32'h00004BBC: begin
				q			<=			16'h2623;
		end
		32'h00004BBE: begin
				q			<=			16'h0CF1;
		end
		32'h00004BC0: begin
				q			<=			16'h2783;
		end
		32'h00004BC2: begin
				q			<=			16'h0C81;
		end
		32'h00004BC4: begin
				q			<=			16'h0713;
		end
		32'h00004BC6: begin
				q			<=			16'h0070;
		end
		32'h00004BC8: begin
				q			<=			16'h8793;
		end
		32'h00004BCA: begin
				q			<=			16'h0017;
		end
		32'h00004BCC: begin
				q			<=			16'h2423;
		end
		32'h00004BCE: begin
				q			<=			16'h0CF1;
		end
		32'h00004BD0: begin
				q			<=			16'h5E63;
		end
		32'h00004BD2: begin
				q			<=			16'h00F7;
		end
		32'h00004BD4: begin
				q			<=			16'h0613;
		end
		32'h00004BD6: begin
				q			<=			16'h0C41;
		end
		32'h00004BD8: begin
				q			<=			16'h8593;
		end
		32'h00004BDA: begin
				q			<=			16'h0009;
		end
		32'h00004BDC: begin
				q			<=			16'h0513;
		end
		32'h00004BDE: begin
				q			<=			16'h0009;
		end
		32'h00004BE0: begin
				q			<=			16'h30EF;
		end
		32'h00004BE2: begin
				q			<=			16'h77D0;
		end
		32'h00004BE4: begin
				q			<=			16'h1663;
		end
		32'h00004BE6: begin
				q			<=			16'h1C05;
		end
		32'h00004BE8: begin
				q			<=			16'h0B93;
		end
		32'h00004BEA: begin
				q			<=			16'h0EC1;
		end
		32'h00004BEC: begin
				q			<=			16'h2783;
		end
		32'h00004BEE: begin
				q			<=			16'h0D01;
		end
		32'h00004BF0: begin
				q			<=			16'h0593;
		end
		32'h00004BF2: begin
				q			<=			16'h0801;
		end
		32'h00004BF4: begin
				q			<=			16'h0513;
		end
		32'h00004BF6: begin
				q			<=			16'h0901;
		end
		32'h00004BF8: begin
				q			<=			16'h2823;
		end
		32'h00004BFA: begin
				q			<=			16'h08F1;
		end
		32'h00004BFC: begin
				q			<=			16'h2783;
		end
		32'h00004BFE: begin
				q			<=			16'h0D41;
		end
		32'h00004C00: begin
				q			<=			16'h0A93;
		end
		32'h00004C02: begin
				q			<=			16'hFFFA;
		end
		32'h00004C04: begin
				q			<=			16'h2023;
		end
		32'h00004C06: begin
				q			<=			16'h0801;
		end
		32'h00004C08: begin
				q			<=			16'h2A23;
		end
		32'h00004C0A: begin
				q			<=			16'h08F1;
		end
		32'h00004C0C: begin
				q			<=			16'h2783;
		end
		32'h00004C0E: begin
				q			<=			16'h0D81;
		end
		32'h00004C10: begin
				q			<=			16'h2223;
		end
		32'h00004C12: begin
				q			<=			16'h0801;
		end
		32'h00004C14: begin
				q			<=			16'h2423;
		end
		32'h00004C16: begin
				q			<=			16'h0801;
		end
		32'h00004C18: begin
				q			<=			16'h2C23;
		end
		32'h00004C1A: begin
				q			<=			16'h08F1;
		end
		32'h00004C1C: begin
				q			<=			16'h2783;
		end
		32'h00004C1E: begin
				q			<=			16'h0DC1;
		end
		32'h00004C20: begin
				q			<=			16'h2623;
		end
		32'h00004C22: begin
				q			<=			16'h0801;
		end
		32'h00004C24: begin
				q			<=			16'h2E23;
		end
		32'h00004C26: begin
				q			<=			16'h08F1;
		end
		32'h00004C28: begin
				q			<=			16'h70EF;
		end
		32'h00004C2A: begin
				q			<=			16'h3940;
		end
		32'h00004C2C: begin
				q			<=			16'h0663;
		end
		32'h00004C2E: begin
				q			<=			16'h0805;
		end
		32'h00004C30: begin
				q			<=			16'h2783;
		end
		32'h00004C32: begin
				q			<=			16'h0CC1;
		end
		32'h00004C34: begin
				q			<=			16'h2703;
		end
		32'h00004C36: begin
				q			<=			16'h0C81;
		end
		32'h00004C38: begin
				q			<=			16'h8493;
		end
		32'h00004C3A: begin
				q			<=			16'h0014;
		end
		32'h00004C3C: begin
				q			<=			16'h8793;
		end
		32'h00004C3E: begin
				q			<=			16'hFFF7;
		end
		32'h00004C40: begin
				q			<=			16'h87B3;
		end
		32'h00004C42: begin
				q			<=			16'h0147;
		end
		32'h00004C44: begin
				q			<=			16'h0713;
		end
		32'h00004C46: begin
				q			<=			16'h0017;
		end
		32'h00004C48: begin
				q			<=			16'hA023;
		end
		32'h00004C4A: begin
				q			<=			16'h009B;
		end
		32'h00004C4C: begin
				q			<=			16'hA223;
		end
		32'h00004C4E: begin
				q			<=			16'h015B;
		end
		32'h00004C50: begin
				q			<=			16'h2623;
		end
		32'h00004C52: begin
				q			<=			16'h0CF1;
		end
		32'h00004C54: begin
				q			<=			16'h2423;
		end
		32'h00004C56: begin
				q			<=			16'h0CE1;
		end
		32'h00004C58: begin
				q			<=			16'h0793;
		end
		32'h00004C5A: begin
				q			<=			16'h0070;
		end
		32'h00004C5C: begin
				q			<=			16'h8B93;
		end
		32'h00004C5E: begin
				q			<=			16'h008B;
		end
		32'h00004C60: begin
				q			<=			16'hDE63;
		end
		32'h00004C62: begin
				q			<=			16'h00E7;
		end
		32'h00004C64: begin
				q			<=			16'h0613;
		end
		32'h00004C66: begin
				q			<=			16'h0C41;
		end
		32'h00004C68: begin
				q			<=			16'h8593;
		end
		32'h00004C6A: begin
				q			<=			16'h0009;
		end
		32'h00004C6C: begin
				q			<=			16'h0513;
		end
		32'h00004C6E: begin
				q			<=			16'h0009;
		end
		32'h00004C70: begin
				q			<=			16'h30EF;
		end
		32'h00004C72: begin
				q			<=			16'h6ED0;
		end
		32'h00004C74: begin
				q			<=			16'h1E63;
		end
		32'h00004C76: begin
				q			<=			16'h1205;
		end
		32'h00004C78: begin
				q			<=			16'h0B93;
		end
		32'h00004C7A: begin
				q			<=			16'h0EC1;
		end
		32'h00004C7C: begin
				q			<=			16'h0793;
		end
		32'h00004C7E: begin
				q			<=			16'h0B41;
		end
		32'h00004C80: begin
				q			<=			16'hA023;
		end
		32'h00004C82: begin
				q			<=			16'h00FB;
		end
		32'h00004C84: begin
				q			<=			16'h2783;
		end
		32'h00004C86: begin
				q			<=			16'h0301;
		end
		32'h00004C88: begin
				q			<=			16'h2703;
		end
		32'h00004C8A: begin
				q			<=			16'h0301;
		end
		32'h00004C8C: begin
				q			<=			16'h8893;
		end
		32'h00004C8E: begin
				q			<=			16'h008B;
		end
		32'h00004C90: begin
				q			<=			16'hA223;
		end
		32'h00004C92: begin
				q			<=			16'h00FB;
		end
		32'h00004C94: begin
				q			<=			16'h2783;
		end
		32'h00004C96: begin
				q			<=			16'h0CC1;
		end
		32'h00004C98: begin
				q			<=			16'h87B3;
		end
		32'h00004C9A: begin
				q			<=			16'h00E7;
		end
		32'h00004C9C: begin
				q			<=			16'h2623;
		end
		32'h00004C9E: begin
				q			<=			16'h0CF1;
		end
		32'h00004CA0: begin
				q			<=			16'h2783;
		end
		32'h00004CA2: begin
				q			<=			16'h0C81;
		end
		32'h00004CA4: begin
				q			<=			16'h0713;
		end
		32'h00004CA6: begin
				q			<=			16'h0070;
		end
		32'h00004CA8: begin
				q			<=			16'h8793;
		end
		32'h00004CAA: begin
				q			<=			16'h0017;
		end
		32'h00004CAC: begin
				q			<=			16'h2423;
		end
		32'h00004CAE: begin
				q			<=			16'h0CF1;
		end
		32'h00004CB0: begin
				q			<=			16'h5AE3;
		end
		32'h00004CB2: begin
				q			<=			16'h8AF7;
		end
		32'h00004CB4: begin
				q			<=			16'hF06F;
		end
		32'h00004CB6: begin
				q			<=			16'hBF0F;
		end
		32'h00004CB8: begin
				q			<=			16'h52E3;
		end
		32'h00004CBA: begin
				q			<=			16'hFD50;
		end
		32'h00004CBC: begin
				q			<=			16'h0C13;
		end
		32'h00004CBE: begin
				q			<=			16'h0100;
		end
		32'h00004CC0: begin
				q			<=			16'hA497;
		end
		32'h00004CC2: begin
				q			<=			16'h0000;
		end
		32'h00004CC4: begin
				q			<=			16'h8493;
		end
		32'h00004CC6: begin
				q			<=			16'h5DC4;
		end
		32'h00004CC8: begin
				q			<=			16'h0D13;
		end
		32'h00004CCA: begin
				q			<=			16'h0070;
		end
		32'h00004CCC: begin
				q			<=			16'h2703;
		end
		32'h00004CCE: begin
				q			<=			16'h0C81;
		end
		32'h00004CD0: begin
				q			<=			16'hA023;
		end
		32'h00004CD2: begin
				q			<=			16'h009B;
		end
		32'h00004CD4: begin
				q			<=			16'h2783;
		end
		32'h00004CD6: begin
				q			<=			16'h0CC1;
		end
		32'h00004CD8: begin
				q			<=			16'h0713;
		end
		32'h00004CDA: begin
				q			<=			16'h0017;
		end
		32'h00004CDC: begin
				q			<=			16'h8693;
		end
		32'h00004CDE: begin
				q			<=			16'h008B;
		end
		32'h00004CE0: begin
				q			<=			16'h4063;
		end
		32'h00004CE2: begin
				q			<=			16'h035C;
		end
		32'h00004CE4: begin
				q			<=			16'h87B3;
		end
		32'h00004CE6: begin
				q			<=			16'h00FA;
		end
		32'h00004CE8: begin
				q			<=			16'hA223;
		end
		32'h00004CEA: begin
				q			<=			16'h015B;
		end
		32'h00004CEC: begin
				q			<=			16'h2623;
		end
		32'h00004CEE: begin
				q			<=			16'h0CF1;
		end
		32'h00004CF0: begin
				q			<=			16'h2423;
		end
		32'h00004CF2: begin
				q			<=			16'h0CE1;
		end
		32'h00004CF4: begin
				q			<=			16'h0793;
		end
		32'h00004CF6: begin
				q			<=			16'h0070;
		end
		32'h00004CF8: begin
				q			<=			16'h8B93;
		end
		32'h00004CFA: begin
				q			<=			16'h0006;
		end
		32'h00004CFC: begin
				q			<=			16'hF06F;
		end
		32'h00004CFE: begin
				q			<=			16'hF65F;
		end
		32'h00004D00: begin
				q			<=			16'h8793;
		end
		32'h00004D02: begin
				q			<=			16'h0107;
		end
		32'h00004D04: begin
				q			<=			16'hA223;
		end
		32'h00004D06: begin
				q			<=			16'h018B;
		end
		32'h00004D08: begin
				q			<=			16'h2623;
		end
		32'h00004D0A: begin
				q			<=			16'h0CF1;
		end
		32'h00004D0C: begin
				q			<=			16'h2423;
		end
		32'h00004D0E: begin
				q			<=			16'h0CE1;
		end
		32'h00004D10: begin
				q			<=			16'h5E63;
		end
		32'h00004D12: begin
				q			<=			16'h00ED;
		end
		32'h00004D14: begin
				q			<=			16'h0613;
		end
		32'h00004D16: begin
				q			<=			16'h0C41;
		end
		32'h00004D18: begin
				q			<=			16'h8593;
		end
		32'h00004D1A: begin
				q			<=			16'h0009;
		end
		32'h00004D1C: begin
				q			<=			16'h0513;
		end
		32'h00004D1E: begin
				q			<=			16'h0009;
		end
		32'h00004D20: begin
				q			<=			16'h30EF;
		end
		32'h00004D22: begin
				q			<=			16'h63D0;
		end
		32'h00004D24: begin
				q			<=			16'h1663;
		end
		32'h00004D26: begin
				q			<=			16'h0805;
		end
		32'h00004D28: begin
				q			<=			16'h0693;
		end
		32'h00004D2A: begin
				q			<=			16'h0EC1;
		end
		32'h00004D2C: begin
				q			<=			16'h8A93;
		end
		32'h00004D2E: begin
				q			<=			16'hFF0A;
		end
		32'h00004D30: begin
				q			<=			16'h8B93;
		end
		32'h00004D32: begin
				q			<=			16'h0006;
		end
		32'h00004D34: begin
				q			<=			16'hF06F;
		end
		32'h00004D36: begin
				q			<=			16'hF99F;
		end
		32'h00004D38: begin
				q			<=			16'hA223;
		end
		32'h00004D3A: begin
				q			<=			16'h00E8;
		end
		32'h00004D3C: begin
				q			<=			16'h2623;
		end
		32'h00004D3E: begin
				q			<=			16'h0DB1;
		end
		32'h00004D40: begin
				q			<=			16'h2423;
		end
		32'h00004D42: begin
				q			<=			16'h0CF1;
		end
		32'h00004D44: begin
				q			<=			16'h0713;
		end
		32'h00004D46: begin
				q			<=			16'h0070;
		end
		32'h00004D48: begin
				q			<=			16'h5AE3;
		end
		32'h00004D4A: begin
				q			<=			16'hF2F7;
		end
		32'h00004D4C: begin
				q			<=			16'hF06F;
		end
		32'h00004D4E: begin
				q			<=			16'hF19F;
		end
		32'h00004D50: begin
				q			<=			16'h2783;
		end
		32'h00004D52: begin
				q			<=			16'h01C1;
		end
		32'h00004D54: begin
				q			<=			16'h2703;
		end
		32'h00004D56: begin
				q			<=			16'h0201;
		end
		32'h00004D58: begin
				q			<=			16'h8433;
		end
		32'h00004D5A: begin
				q			<=			16'h40E7;
		end
		32'h00004D5C: begin
				q			<=			16'h58E3;
		end
		32'h00004D5E: begin
				q			<=			16'h8080;
		end
		32'h00004D60: begin
				q			<=			16'h0A93;
		end
		32'h00004D62: begin
				q			<=			16'h0100;
		end
		32'h00004D64: begin
				q			<=			16'hA497;
		end
		32'h00004D66: begin
				q			<=			16'h0000;
		end
		32'h00004D68: begin
				q			<=			16'h8493;
		end
		32'h00004D6A: begin
				q			<=			16'h5284;
		end
		32'h00004D6C: begin
				q			<=			16'h0B93;
		end
		32'h00004D6E: begin
				q			<=			16'h0070;
		end
		32'h00004D70: begin
				q			<=			16'h2783;
		end
		32'h00004D72: begin
				q			<=			16'h0C81;
		end
		32'h00004D74: begin
				q			<=			16'hA023;
		end
		32'h00004D76: begin
				q			<=			16'h0098;
		end
		32'h00004D78: begin
				q			<=			16'h2703;
		end
		32'h00004D7A: begin
				q			<=			16'h0CC1;
		end
		32'h00004D7C: begin
				q			<=			16'h8793;
		end
		32'h00004D7E: begin
				q			<=			16'h0017;
		end
		32'h00004D80: begin
				q			<=			16'hC863;
		end
		32'h00004D82: begin
				q			<=			16'h048A;
		end
		32'h00004D84: begin
				q			<=			16'hA223;
		end
		32'h00004D86: begin
				q			<=			16'h0088;
		end
		32'h00004D88: begin
				q			<=			16'h0433;
		end
		32'h00004D8A: begin
				q			<=			16'h00E4;
		end
		32'h00004D8C: begin
				q			<=			16'h2623;
		end
		32'h00004D8E: begin
				q			<=			16'h0C81;
		end
		32'h00004D90: begin
				q			<=			16'h2423;
		end
		32'h00004D92: begin
				q			<=			16'h0CF1;
		end
		32'h00004D94: begin
				q			<=			16'h0713;
		end
		32'h00004D96: begin
				q			<=			16'h0070;
		end
		32'h00004D98: begin
				q			<=			16'h5A63;
		end
		32'h00004D9A: begin
				q			<=			16'hFCF7;
		end
		32'h00004D9C: begin
				q			<=			16'h0613;
		end
		32'h00004D9E: begin
				q			<=			16'h0C41;
		end
		32'h00004DA0: begin
				q			<=			16'h8593;
		end
		32'h00004DA2: begin
				q			<=			16'h0009;
		end
		32'h00004DA4: begin
				q			<=			16'h0513;
		end
		32'h00004DA6: begin
				q			<=			16'h0009;
		end
		32'h00004DA8: begin
				q			<=			16'h30EF;
		end
		32'h00004DAA: begin
				q			<=			16'h5B50;
		end
		32'h00004DAC: begin
				q			<=			16'h0063;
		end
		32'h00004DAE: begin
				q			<=			16'hFC05;
		end
		32'h00004DB0: begin
				q			<=			16'h2783;
		end
		32'h00004DB2: begin
				q			<=			16'h0041;
		end
		32'h00004DB4: begin
				q			<=			16'h9463;
		end
		32'h00004DB6: begin
				q			<=			16'h0007;
		end
		32'h00004DB8: begin
				q			<=			16'hE06F;
		end
		32'h00004DBA: begin
				q			<=			16'hF48F;
		end
		32'h00004DBC: begin
				q			<=			16'h8593;
		end
		32'h00004DBE: begin
				q			<=			16'h0007;
		end
		32'h00004DC0: begin
				q			<=			16'h0513;
		end
		32'h00004DC2: begin
				q			<=			16'h0009;
		end
		32'h00004DC4: begin
				q			<=			16'h0097;
		end
		32'h00004DC6: begin
				q			<=			16'h0000;
		end
		32'h00004DC8: begin
				q			<=			16'h80E7;
		end
		32'h00004DCA: begin
				q			<=			16'h1AC0;
		end
		32'h00004DCC: begin
				q			<=			16'hE06F;
		end
		32'h00004DCE: begin
				q			<=			16'hF34F;
		end
		32'h00004DD0: begin
				q			<=			16'h0713;
		end
		32'h00004DD2: begin
				q			<=			16'h0107;
		end
		32'h00004DD4: begin
				q			<=			16'hA223;
		end
		32'h00004DD6: begin
				q			<=			16'h0158;
		end
		32'h00004DD8: begin
				q			<=			16'h2623;
		end
		32'h00004DDA: begin
				q			<=			16'h0CE1;
		end
		32'h00004DDC: begin
				q			<=			16'h2423;
		end
		32'h00004DDE: begin
				q			<=			16'h0CF1;
		end
		32'h00004DE0: begin
				q			<=			16'h8893;
		end
		32'h00004DE2: begin
				q			<=			16'h0088;
		end
		32'h00004DE4: begin
				q			<=			16'hDE63;
		end
		32'h00004DE6: begin
				q			<=			16'h00FB;
		end
		32'h00004DE8: begin
				q			<=			16'h0613;
		end
		32'h00004DEA: begin
				q			<=			16'h0C41;
		end
		32'h00004DEC: begin
				q			<=			16'h8593;
		end
		32'h00004DEE: begin
				q			<=			16'h0009;
		end
		32'h00004DF0: begin
				q			<=			16'h0513;
		end
		32'h00004DF2: begin
				q			<=			16'h0009;
		end
		32'h00004DF4: begin
				q			<=			16'h30EF;
		end
		32'h00004DF6: begin
				q			<=			16'h5690;
		end
		32'h00004DF8: begin
				q			<=			16'h1CE3;
		end
		32'h00004DFA: begin
				q			<=			16'hFA05;
		end
		32'h00004DFC: begin
				q			<=			16'h0893;
		end
		32'h00004DFE: begin
				q			<=			16'h0EC1;
		end
		32'h00004E00: begin
				q			<=			16'h0413;
		end
		32'h00004E02: begin
				q			<=			16'hFF04;
		end
		32'h00004E04: begin
				q			<=			16'hF06F;
		end
		32'h00004E06: begin
				q			<=			16'hF6DF;
		end
		32'h00004E08: begin
				q			<=			16'h2583;
		end
		32'h00004E0A: begin
				q			<=			16'h0041;
		end
		32'h00004E0C: begin
				q			<=			16'h0513;
		end
		32'h00004E0E: begin
				q			<=			16'h0009;
		end
		32'h00004E10: begin
				q			<=			16'h0097;
		end
		32'h00004E12: begin
				q			<=			16'h0000;
		end
		32'h00004E14: begin
				q			<=			16'h80E7;
		end
		32'h00004E16: begin
				q			<=			16'h1600;
		end
		32'h00004E18: begin
				q			<=			16'hF06F;
		end
		32'h00004E1A: begin
				q			<=			16'hF98F;
		end
		32'h00004E1C: begin
				q			<=			16'h2783;
		end
		32'h00004E1E: begin
				q			<=			16'h0CC1;
		end
		32'h00004E20: begin
				q			<=			16'h9463;
		end
		32'h00004E22: begin
				q			<=			16'h0007;
		end
		32'h00004E24: begin
				q			<=			16'hE06F;
		end
		32'h00004E26: begin
				q			<=			16'hEDCF;
		end
		32'h00004E28: begin
				q			<=			16'h0613;
		end
		32'h00004E2A: begin
				q			<=			16'h0C41;
		end
		32'h00004E2C: begin
				q			<=			16'h8593;
		end
		32'h00004E2E: begin
				q			<=			16'h0009;
		end
		32'h00004E30: begin
				q			<=			16'h0513;
		end
		32'h00004E32: begin
				q			<=			16'h0009;
		end
		32'h00004E34: begin
				q			<=			16'h30EF;
		end
		32'h00004E36: begin
				q			<=			16'h5290;
		end
		32'h00004E38: begin
				q			<=			16'hE06F;
		end
		32'h00004E3A: begin
				q			<=			16'hEC8F;
		end
		32'h00004E3C: begin
				q			<=			16'h0000;
		end
		32'h00004E3E: begin
				q			<=			16'h0000;
		end
		32'h00004E40: begin
				q			<=			16'h0113;
		end
		32'h00004E42: begin
				q			<=			16'hFD01;
		end
		32'h00004E44: begin
				q			<=			16'h2423;
		end
		32'h00004E46: begin
				q			<=			16'h0281;
		end
		32'h00004E48: begin
				q			<=			16'h2223;
		end
		32'h00004E4A: begin
				q			<=			16'h0291;
		end
		32'h00004E4C: begin
				q			<=			16'h2023;
		end
		32'h00004E4E: begin
				q			<=			16'h0321;
		end
		32'h00004E50: begin
				q			<=			16'h2E23;
		end
		32'h00004E52: begin
				q			<=			16'h0131;
		end
		32'h00004E54: begin
				q			<=			16'h2623;
		end
		32'h00004E56: begin
				q			<=			16'h00B1;
		end
		32'h00004E58: begin
				q			<=			16'h2623;
		end
		32'h00004E5A: begin
				q			<=			16'h0211;
		end
		32'h00004E5C: begin
				q			<=			16'h0913;
		end
		32'h00004E5E: begin
				q			<=			16'h0005;
		end
		32'h00004E60: begin
				q			<=			16'hB997;
		end
		32'h00004E62: begin
				q			<=			16'h0000;
		end
		32'h00004E64: begin
				q			<=			16'h8993;
		end
		32'h00004E66: begin
				q			<=			16'h5009;
		end
		32'h00004E68: begin
				q			<=			16'h20EF;
		end
		32'h00004E6A: begin
				q			<=			16'h4190;
		end
		32'h00004E6C: begin
				q			<=			16'hA783;
		end
		32'h00004E6E: begin
				q			<=			16'h0089;
		end
		32'h00004E70: begin
				q			<=			16'h2583;
		end
		32'h00004E72: begin
				q			<=			16'h00C1;
		end
		32'h00004E74: begin
				q			<=			16'hA483;
		end
		32'h00004E76: begin
				q			<=			16'h0047;
		end
		32'h00004E78: begin
				q			<=			16'h17B7;
		end
		32'h00004E7A: begin
				q			<=			16'h0000;
		end
		32'h00004E7C: begin
				q			<=			16'h8413;
		end
		32'h00004E7E: begin
				q			<=			16'hFEF7;
		end
		32'h00004E80: begin
				q			<=			16'hF493;
		end
		32'h00004E82: begin
				q			<=			16'hFFC4;
		end
		32'h00004E84: begin
				q			<=			16'h0433;
		end
		32'h00004E86: begin
				q			<=			16'h40B4;
		end
		32'h00004E88: begin
				q			<=			16'h0433;
		end
		32'h00004E8A: begin
				q			<=			16'h0094;
		end
		32'h00004E8C: begin
				q			<=			16'h5413;
		end
		32'h00004E8E: begin
				q			<=			16'h00C4;
		end
		32'h00004E90: begin
				q			<=			16'h0413;
		end
		32'h00004E92: begin
				q			<=			16'hFFF4;
		end
		32'h00004E94: begin
				q			<=			16'h1413;
		end
		32'h00004E96: begin
				q			<=			16'h00C4;
		end
		32'h00004E98: begin
				q			<=			16'h5863;
		end
		32'h00004E9A: begin
				q			<=			16'h02F4;
		end
		32'h00004E9C: begin
				q			<=			16'h0513;
		end
		32'h00004E9E: begin
				q			<=			16'h0009;
		end
		32'h00004EA0: begin
				q			<=			16'h3097;
		end
		32'h00004EA2: begin
				q			<=			16'h0000;
		end
		32'h00004EA4: begin
				q			<=			16'h80E7;
		end
		32'h00004EA6: begin
				q			<=			16'hBE40;
		end
		32'h00004EA8: begin
				q			<=			16'h0513;
		end
		32'h00004EAA: begin
				q			<=			16'h0000;
		end
		32'h00004EAC: begin
				q			<=			16'h2083;
		end
		32'h00004EAE: begin
				q			<=			16'h02C1;
		end
		32'h00004EB0: begin
				q			<=			16'h2403;
		end
		32'h00004EB2: begin
				q			<=			16'h0281;
		end
		32'h00004EB4: begin
				q			<=			16'h2483;
		end
		32'h00004EB6: begin
				q			<=			16'h0241;
		end
		32'h00004EB8: begin
				q			<=			16'h2903;
		end
		32'h00004EBA: begin
				q			<=			16'h0201;
		end
		32'h00004EBC: begin
				q			<=			16'h2983;
		end
		32'h00004EBE: begin
				q			<=			16'h01C1;
		end
		32'h00004EC0: begin
				q			<=			16'h0113;
		end
		32'h00004EC2: begin
				q			<=			16'h0301;
		end
		32'h00004EC4: begin
				q			<=			16'h8067;
		end
		32'h00004EC6: begin
				q			<=			16'h0000;
		end
		32'h00004EC8: begin
				q			<=			16'h0593;
		end
		32'h00004ECA: begin
				q			<=			16'h0000;
		end
		32'h00004ECC: begin
				q			<=			16'h0513;
		end
		32'h00004ECE: begin
				q			<=			16'h0009;
		end
		32'h00004ED0: begin
				q			<=			16'h30EF;
		end
		32'h00004ED2: begin
				q			<=			16'h3390;
		end
		32'h00004ED4: begin
				q			<=			16'hA783;
		end
		32'h00004ED6: begin
				q			<=			16'h0089;
		end
		32'h00004ED8: begin
				q			<=			16'h87B3;
		end
		32'h00004EDA: begin
				q			<=			16'h0097;
		end
		32'h00004EDC: begin
				q			<=			16'h10E3;
		end
		32'h00004EDE: begin
				q			<=			16'hFCF5;
		end
		32'h00004EE0: begin
				q			<=			16'h05B3;
		end
		32'h00004EE2: begin
				q			<=			16'h4080;
		end
		32'h00004EE4: begin
				q			<=			16'h0513;
		end
		32'h00004EE6: begin
				q			<=			16'h0009;
		end
		32'h00004EE8: begin
				q			<=			16'h30EF;
		end
		32'h00004EEA: begin
				q			<=			16'h3210;
		end
		32'h00004EEC: begin
				q			<=			16'h0793;
		end
		32'h00004EEE: begin
				q			<=			16'hFFF0;
		end
		32'h00004EF0: begin
				q			<=			16'h1263;
		end
		32'h00004EF2: begin
				q			<=			16'h04F5;
		end
		32'h00004EF4: begin
				q			<=			16'h0593;
		end
		32'h00004EF6: begin
				q			<=			16'h0000;
		end
		32'h00004EF8: begin
				q			<=			16'h0513;
		end
		32'h00004EFA: begin
				q			<=			16'h0009;
		end
		32'h00004EFC: begin
				q			<=			16'h30EF;
		end
		32'h00004EFE: begin
				q			<=			16'h30D0;
		end
		32'h00004F00: begin
				q			<=			16'hA703;
		end
		32'h00004F02: begin
				q			<=			16'h0089;
		end
		32'h00004F04: begin
				q			<=			16'h0693;
		end
		32'h00004F06: begin
				q			<=			16'h00F0;
		end
		32'h00004F08: begin
				q			<=			16'h07B3;
		end
		32'h00004F0A: begin
				q			<=			16'h40E5;
		end
		32'h00004F0C: begin
				q			<=			16'hD8E3;
		end
		32'h00004F0E: begin
				q			<=			16'hF8F6;
		end
		32'h00004F10: begin
				q			<=			16'hC697;
		end
		32'h00004F12: begin
				q			<=			16'h0000;
		end
		32'h00004F14: begin
				q			<=			16'h8693;
		end
		32'h00004F16: begin
				q			<=			16'h9CC6;
		end
		32'h00004F18: begin
				q			<=			16'hA683;
		end
		32'h00004F1A: begin
				q			<=			16'h0006;
		end
		32'h00004F1C: begin
				q			<=			16'hE793;
		end
		32'h00004F1E: begin
				q			<=			16'h0017;
		end
		32'h00004F20: begin
				q			<=			16'h2223;
		end
		32'h00004F22: begin
				q			<=			16'h00F7;
		end
		32'h00004F24: begin
				q			<=			16'h0533;
		end
		32'h00004F26: begin
				q			<=			16'h40D5;
		end
		32'h00004F28: begin
				q			<=			16'hC697;
		end
		32'h00004F2A: begin
				q			<=			16'h0000;
		end
		32'h00004F2C: begin
				q			<=			16'hA623;
		end
		32'h00004F2E: begin
				q			<=			16'hBCA6;
		end
		32'h00004F30: begin
				q			<=			16'hF06F;
		end
		32'h00004F32: begin
				q			<=			16'hF6DF;
		end
		32'h00004F34: begin
				q			<=			16'hA783;
		end
		32'h00004F36: begin
				q			<=			16'h0089;
		end
		32'h00004F38: begin
				q			<=			16'h84B3;
		end
		32'h00004F3A: begin
				q			<=			16'h4084;
		end
		32'h00004F3C: begin
				q			<=			16'hE493;
		end
		32'h00004F3E: begin
				q			<=			16'h0014;
		end
		32'h00004F40: begin
				q			<=			16'hA223;
		end
		32'h00004F42: begin
				q			<=			16'h0097;
		end
		32'h00004F44: begin
				q			<=			16'hC797;
		end
		32'h00004F46: begin
				q			<=			16'h0000;
		end
		32'h00004F48: begin
				q			<=			16'h8793;
		end
		32'h00004F4A: begin
				q			<=			16'hBB07;
		end
		32'h00004F4C: begin
				q			<=			16'hA783;
		end
		32'h00004F4E: begin
				q			<=			16'h0007;
		end
		32'h00004F50: begin
				q			<=			16'h0513;
		end
		32'h00004F52: begin
				q			<=			16'h0009;
		end
		32'h00004F54: begin
				q			<=			16'h8433;
		end
		32'h00004F56: begin
				q			<=			16'h4087;
		end
		32'h00004F58: begin
				q			<=			16'hC797;
		end
		32'h00004F5A: begin
				q			<=			16'h0000;
		end
		32'h00004F5C: begin
				q			<=			16'hAE23;
		end
		32'h00004F5E: begin
				q			<=			16'hB887;
		end
		32'h00004F60: begin
				q			<=			16'h3097;
		end
		32'h00004F62: begin
				q			<=			16'h0000;
		end
		32'h00004F64: begin
				q			<=			16'h80E7;
		end
		32'h00004F66: begin
				q			<=			16'hB240;
		end
		32'h00004F68: begin
				q			<=			16'h0513;
		end
		32'h00004F6A: begin
				q			<=			16'h0010;
		end
		32'h00004F6C: begin
				q			<=			16'hF06F;
		end
		32'h00004F6E: begin
				q			<=			16'hF41F;
		end
		32'h00004F70: begin
				q			<=			16'h8063;
		end
		32'h00004F72: begin
				q			<=			16'h2805;
		end
		32'h00004F74: begin
				q			<=			16'h0113;
		end
		32'h00004F76: begin
				q			<=			16'hFF01;
		end
		32'h00004F78: begin
				q			<=			16'h2423;
		end
		32'h00004F7A: begin
				q			<=			16'h0081;
		end
		32'h00004F7C: begin
				q			<=			16'h2223;
		end
		32'h00004F7E: begin
				q			<=			16'h0091;
		end
		32'h00004F80: begin
				q			<=			16'h0413;
		end
		32'h00004F82: begin
				q			<=			16'h0005;
		end
		32'h00004F84: begin
				q			<=			16'h8493;
		end
		32'h00004F86: begin
				q			<=			16'h0005;
		end
		32'h00004F88: begin
				q			<=			16'h2623;
		end
		32'h00004F8A: begin
				q			<=			16'h0011;
		end
		32'h00004F8C: begin
				q			<=			16'h3097;
		end
		32'h00004F8E: begin
				q			<=			16'h0000;
		end
		32'h00004F90: begin
				q			<=			16'h80E7;
		end
		32'h00004F92: begin
				q			<=			16'hAF40;
		end
		32'h00004F94: begin
				q			<=			16'hA583;
		end
		32'h00004F96: begin
				q			<=			16'hFFC4;
		end
		32'h00004F98: begin
				q			<=			16'h8693;
		end
		32'h00004F9A: begin
				q			<=			16'hFF84;
		end
		32'h00004F9C: begin
				q			<=			16'hB517;
		end
		32'h00004F9E: begin
				q			<=			16'h0000;
		end
		32'h00004FA0: begin
				q			<=			16'h0513;
		end
		32'h00004FA2: begin
				q			<=			16'h3C45;
		end
		32'h00004FA4: begin
				q			<=			16'hF793;
		end
		32'h00004FA6: begin
				q			<=			16'hFFE5;
		end
		32'h00004FA8: begin
				q			<=			16'h8633;
		end
		32'h00004FAA: begin
				q			<=			16'h00F6;
		end
		32'h00004FAC: begin
				q			<=			16'h2703;
		end
		32'h00004FAE: begin
				q			<=			16'h0046;
		end
		32'h00004FB0: begin
				q			<=			16'h2803;
		end
		32'h00004FB2: begin
				q			<=			16'h0085;
		end
		32'h00004FB4: begin
				q			<=			16'hF593;
		end
		32'h00004FB6: begin
				q			<=			16'h0015;
		end
		32'h00004FB8: begin
				q			<=			16'h7713;
		end
		32'h00004FBA: begin
				q			<=			16'hFFC7;
		end
		32'h00004FBC: begin
				q			<=			16'h1C63;
		end
		32'h00004FBE: begin
				q			<=			16'h06C8;
		end
		32'h00004FC0: begin
				q			<=			16'h87B3;
		end
		32'h00004FC2: begin
				q			<=			16'h00E7;
		end
		32'h00004FC4: begin
				q			<=			16'h9063;
		end
		32'h00004FC6: begin
				q			<=			16'h0205;
		end
		32'h00004FC8: begin
				q			<=			16'hA703;
		end
		32'h00004FCA: begin
				q			<=			16'hFF84;
		end
		32'h00004FCC: begin
				q			<=			16'h86B3;
		end
		32'h00004FCE: begin
				q			<=			16'h40E6;
		end
		32'h00004FD0: begin
				q			<=			16'hA603;
		end
		32'h00004FD2: begin
				q			<=			16'h0086;
		end
		32'h00004FD4: begin
				q			<=			16'h87B3;
		end
		32'h00004FD6: begin
				q			<=			16'h00E7;
		end
		32'h00004FD8: begin
				q			<=			16'hA703;
		end
		32'h00004FDA: begin
				q			<=			16'h00C6;
		end
		32'h00004FDC: begin
				q			<=			16'h2623;
		end
		32'h00004FDE: begin
				q			<=			16'h00E6;
		end
		32'h00004FE0: begin
				q			<=			16'h2423;
		end
		32'h00004FE2: begin
				q			<=			16'h00C7;
		end
		32'h00004FE4: begin
				q			<=			16'hE713;
		end
		32'h00004FE6: begin
				q			<=			16'h0017;
		end
		32'h00004FE8: begin
				q			<=			16'hA223;
		end
		32'h00004FEA: begin
				q			<=			16'h00E6;
		end
		32'h00004FEC: begin
				q			<=			16'hB717;
		end
		32'h00004FEE: begin
				q			<=			16'h0000;
		end
		32'h00004FF0: begin
				q			<=			16'h2E23;
		end
		32'h00004FF2: begin
				q			<=			16'h36D7;
		end
		32'h00004FF4: begin
				q			<=			16'hC717;
		end
		32'h00004FF6: begin
				q			<=			16'h0000;
		end
		32'h00004FF8: begin
				q			<=			16'h0713;
		end
		32'h00004FFA: begin
				q			<=			16'h8EC7;
		end
		32'h00004FFC: begin
				q			<=			16'h2703;
		end
		32'h00004FFE: begin
				q			<=			16'h0007;
		end
		32'h00005000: begin
				q			<=			16'hEE63;
		end
		32'h00005002: begin
				q			<=			16'h00E7;
		end
		32'h00005004: begin
				q			<=			16'hC797;
		end
		32'h00005006: begin
				q			<=			16'h0000;
		end
		32'h00005008: begin
				q			<=			16'h8793;
		end
		32'h0000500A: begin
				q			<=			16'hFA47;
		end
		32'h0000500C: begin
				q			<=			16'hA583;
		end
		32'h0000500E: begin
				q			<=			16'h0007;
		end
		32'h00005010: begin
				q			<=			16'h0513;
		end
		32'h00005012: begin
				q			<=			16'h0004;
		end
		32'h00005014: begin
				q			<=			16'h0097;
		end
		32'h00005016: begin
				q			<=			16'h0000;
		end
		32'h00005018: begin
				q			<=			16'h80E7;
		end
		32'h0000501A: begin
				q			<=			16'hE2C0;
		end
		32'h0000501C: begin
				q			<=			16'h0513;
		end
		32'h0000501E: begin
				q			<=			16'h0004;
		end
		32'h00005020: begin
				q			<=			16'h2403;
		end
		32'h00005022: begin
				q			<=			16'h0081;
		end
		32'h00005024: begin
				q			<=			16'h2083;
		end
		32'h00005026: begin
				q			<=			16'h00C1;
		end
		32'h00005028: begin
				q			<=			16'h2483;
		end
		32'h0000502A: begin
				q			<=			16'h0041;
		end
		32'h0000502C: begin
				q			<=			16'h0113;
		end
		32'h0000502E: begin
				q			<=			16'h0101;
		end
		32'h00005030: begin
				q			<=			16'h206F;
		end
		32'h00005032: begin
				q			<=			16'h2550;
		end
		32'h00005034: begin
				q			<=			16'h2223;
		end
		32'h00005036: begin
				q			<=			16'h00E6;
		end
		32'h00005038: begin
				q			<=			16'h0813;
		end
		32'h0000503A: begin
				q			<=			16'h0000;
		end
		32'h0000503C: begin
				q			<=			16'h9663;
		end
		32'h0000503E: begin
				q			<=			16'h0205;
		end
		32'h00005040: begin
				q			<=			16'hA583;
		end
		32'h00005042: begin
				q			<=			16'hFF84;
		end
		32'h00005044: begin
				q			<=			16'hB897;
		end
		32'h00005046: begin
				q			<=			16'h0000;
		end
		32'h00005048: begin
				q			<=			16'h8893;
		end
		32'h0000504A: begin
				q			<=			16'h3248;
		end
		32'h0000504C: begin
				q			<=			16'h86B3;
		end
		32'h0000504E: begin
				q			<=			16'h40B6;
		end
		32'h00005050: begin
				q			<=			16'h87B3;
		end
		32'h00005052: begin
				q			<=			16'h00B7;
		end
		32'h00005054: begin
				q			<=			16'hA583;
		end
		32'h00005056: begin
				q			<=			16'h0086;
		end
		32'h00005058: begin
				q			<=			16'h8C63;
		end
		32'h0000505A: begin
				q			<=			16'h0B15;
		end
		32'h0000505C: begin
				q			<=			16'hA883;
		end
		32'h0000505E: begin
				q			<=			16'h00C6;
		end
		32'h00005060: begin
				q			<=			16'hA623;
		end
		32'h00005062: begin
				q			<=			16'h0115;
		end
		32'h00005064: begin
				q			<=			16'hA423;
		end
		32'h00005066: begin
				q			<=			16'h00B8;
		end
		32'h00005068: begin
				q			<=			16'h05B3;
		end
		32'h0000506A: begin
				q			<=			16'h00E6;
		end
		32'h0000506C: begin
				q			<=			16'hA583;
		end
		32'h0000506E: begin
				q			<=			16'h0045;
		end
		32'h00005070: begin
				q			<=			16'hF593;
		end
		32'h00005072: begin
				q			<=			16'h0015;
		end
		32'h00005074: begin
				q			<=			16'h9C63;
		end
		32'h00005076: begin
				q			<=			16'h0205;
		end
		32'h00005078: begin
				q			<=			16'h87B3;
		end
		32'h0000507A: begin
				q			<=			16'h00E7;
		end
		32'h0000507C: begin
				q			<=			16'h2703;
		end
		32'h0000507E: begin
				q			<=			16'h0086;
		end
		32'h00005080: begin
				q			<=			16'h1C63;
		end
		32'h00005082: begin
				q			<=			16'h0808;
		end
		32'h00005084: begin
				q			<=			16'hB597;
		end
		32'h00005086: begin
				q			<=			16'h0000;
		end
		32'h00005088: begin
				q			<=			16'h8593;
		end
		32'h0000508A: begin
				q			<=			16'h2E45;
		end
		32'h0000508C: begin
				q			<=			16'h1663;
		end
		32'h0000508E: begin
				q			<=			16'h08B7;
		end
		32'h00005090: begin
				q			<=			16'hB617;
		end
		32'h00005092: begin
				q			<=			16'h0000;
		end
		32'h00005094: begin
				q			<=			16'h2223;
		end
		32'h00005096: begin
				q			<=			16'h2ED6;
		end
		32'h00005098: begin
				q			<=			16'hB617;
		end
		32'h0000509A: begin
				q			<=			16'h0000;
		end
		32'h0000509C: begin
				q			<=			16'h2C23;
		end
		32'h0000509E: begin
				q			<=			16'h2CD6;
		end
		32'h000050A0: begin
				q			<=			16'hA623;
		end
		32'h000050A2: begin
				q			<=			16'h00E6;
		end
		32'h000050A4: begin
				q			<=			16'hA423;
		end
		32'h000050A6: begin
				q			<=			16'h00E6;
		end
		32'h000050A8: begin
				q			<=			16'h0813;
		end
		32'h000050AA: begin
				q			<=			16'h0010;
		end
		32'h000050AC: begin
				q			<=			16'hE713;
		end
		32'h000050AE: begin
				q			<=			16'h0017;
		end
		32'h000050B0: begin
				q			<=			16'hA223;
		end
		32'h000050B2: begin
				q			<=			16'h00E6;
		end
		32'h000050B4: begin
				q			<=			16'h8733;
		end
		32'h000050B6: begin
				q			<=			16'h00F6;
		end
		32'h000050B8: begin
				q			<=			16'h2023;
		end
		32'h000050BA: begin
				q			<=			16'h00F7;
		end
		32'h000050BC: begin
				q			<=			16'h10E3;
		end
		32'h000050BE: begin
				q			<=			16'hF608;
		end
		32'h000050C0: begin
				q			<=			16'h0713;
		end
		32'h000050C2: begin
				q			<=			16'h1FF0;
		end
		32'h000050C4: begin
				q			<=			16'h6263;
		end
		32'h000050C6: begin
				q			<=			16'h06F7;
		end
		32'h000050C8: begin
				q			<=			16'hD793;
		end
		32'h000050CA: begin
				q			<=			16'h0037;
		end
		32'h000050CC: begin
				q			<=			16'hD613;
		end
		32'h000050CE: begin
				q			<=			16'h4027;
		end
		32'h000050D0: begin
				q			<=			16'h0713;
		end
		32'h000050D2: begin
				q			<=			16'h0010;
		end
		32'h000050D4: begin
				q			<=			16'h1733;
		end
		32'h000050D6: begin
				q			<=			16'h00C7;
		end
		32'h000050D8: begin
				q			<=			16'h2603;
		end
		32'h000050DA: begin
				q			<=			16'h0045;
		end
		32'h000050DC: begin
				q			<=			16'h8793;
		end
		32'h000050DE: begin
				q			<=			16'h0017;
		end
		32'h000050E0: begin
				q			<=			16'h9793;
		end
		32'h000050E2: begin
				q			<=			16'h0037;
		end
		32'h000050E4: begin
				q			<=			16'h6733;
		end
		32'h000050E6: begin
				q			<=			16'h00C7;
		end
		32'h000050E8: begin
				q			<=			16'h07B3;
		end
		32'h000050EA: begin
				q			<=			16'h00F5;
		end
		32'h000050EC: begin
				q			<=			16'hB617;
		end
		32'h000050EE: begin
				q			<=			16'h0000;
		end
		32'h000050F0: begin
				q			<=			16'h2C23;
		end
		32'h000050F2: begin
				q			<=			16'h26E6;
		end
		32'h000050F4: begin
				q			<=			16'hA703;
		end
		32'h000050F6: begin
				q			<=			16'h0007;
		end
		32'h000050F8: begin
				q			<=			16'h8613;
		end
		32'h000050FA: begin
				q			<=			16'hFF87;
		end
		32'h000050FC: begin
				q			<=			16'hA623;
		end
		32'h000050FE: begin
				q			<=			16'h00C6;
		end
		32'h00005100: begin
				q			<=			16'hA423;
		end
		32'h00005102: begin
				q			<=			16'h00E6;
		end
		32'h00005104: begin
				q			<=			16'hA023;
		end
		32'h00005106: begin
				q			<=			16'h00D7;
		end
		32'h00005108: begin
				q			<=			16'h2623;
		end
		32'h0000510A: begin
				q			<=			16'h00D7;
		end
		32'h0000510C: begin
				q			<=			16'hF06F;
		end
		32'h0000510E: begin
				q			<=			16'hF11F;
		end
		32'h00005110: begin
				q			<=			16'h0813;
		end
		32'h00005112: begin
				q			<=			16'h0010;
		end
		32'h00005114: begin
				q			<=			16'hF06F;
		end
		32'h00005116: begin
				q			<=			16'hF55F;
		end
		32'h00005118: begin
				q			<=			16'h2603;
		end
		32'h0000511A: begin
				q			<=			16'h00C6;
		end
		32'h0000511C: begin
				q			<=			16'h2623;
		end
		32'h0000511E: begin
				q			<=			16'h00C7;
		end
		32'h00005120: begin
				q			<=			16'h2423;
		end
		32'h00005122: begin
				q			<=			16'h00E6;
		end
		32'h00005124: begin
				q			<=			16'hF06F;
		end
		32'h00005126: begin
				q			<=			16'hF89F;
		end
		32'h00005128: begin
				q			<=			16'hD613;
		end
		32'h0000512A: begin
				q			<=			16'h0097;
		end
		32'h0000512C: begin
				q			<=			16'h0713;
		end
		32'h0000512E: begin
				q			<=			16'h0040;
		end
		32'h00005130: begin
				q			<=			16'h6A63;
		end
		32'h00005132: begin
				q			<=			16'h04C7;
		end
		32'h00005134: begin
				q			<=			16'hD713;
		end
		32'h00005136: begin
				q			<=			16'h0067;
		end
		32'h00005138: begin
				q			<=			16'h0713;
		end
		32'h0000513A: begin
				q			<=			16'h0387;
		end
		32'h0000513C: begin
				q			<=			16'h0613;
		end
		32'h0000513E: begin
				q			<=			16'h0017;
		end
		32'h00005140: begin
				q			<=			16'h1613;
		end
		32'h00005142: begin
				q			<=			16'h0036;
		end
		32'h00005144: begin
				q			<=			16'h0633;
		end
		32'h00005146: begin
				q			<=			16'h00C5;
		end
		32'h00005148: begin
				q			<=			16'h0593;
		end
		32'h0000514A: begin
				q			<=			16'hFF86;
		end
		32'h0000514C: begin
				q			<=			16'h2603;
		end
		32'h0000514E: begin
				q			<=			16'h0006;
		end
		32'h00005150: begin
				q			<=			16'h9663;
		end
		32'h00005152: begin
				q			<=			16'h08C5;
		end
		32'h00005154: begin
				q			<=			16'h0793;
		end
		32'h00005156: begin
				q			<=			16'h0010;
		end
		32'h00005158: begin
				q			<=			16'h5713;
		end
		32'h0000515A: begin
				q			<=			16'h4027;
		end
		32'h0000515C: begin
				q			<=			16'h9733;
		end
		32'h0000515E: begin
				q			<=			16'h00E7;
		end
		32'h00005160: begin
				q			<=			16'h2783;
		end
		32'h00005162: begin
				q			<=			16'h0045;
		end
		32'h00005164: begin
				q			<=			16'h6733;
		end
		32'h00005166: begin
				q			<=			16'h00F7;
		end
		32'h00005168: begin
				q			<=			16'hB797;
		end
		32'h0000516A: begin
				q			<=			16'h0000;
		end
		32'h0000516C: begin
				q			<=			16'hAE23;
		end
		32'h0000516E: begin
				q			<=			16'h1EE7;
		end
		32'h00005170: begin
				q			<=			16'hA623;
		end
		32'h00005172: begin
				q			<=			16'h00B6;
		end
		32'h00005174: begin
				q			<=			16'hA423;
		end
		32'h00005176: begin
				q			<=			16'h00C6;
		end
		32'h00005178: begin
				q			<=			16'hA423;
		end
		32'h0000517A: begin
				q			<=			16'h00D5;
		end
		32'h0000517C: begin
				q			<=			16'h2623;
		end
		32'h0000517E: begin
				q			<=			16'h00D6;
		end
		32'h00005180: begin
				q			<=			16'hF06F;
		end
		32'h00005182: begin
				q			<=			16'hE9DF;
		end
		32'h00005184: begin
				q			<=			16'h0713;
		end
		32'h00005186: begin
				q			<=			16'h0140;
		end
		32'h00005188: begin
				q			<=			16'h6663;
		end
		32'h0000518A: begin
				q			<=			16'h00C7;
		end
		32'h0000518C: begin
				q			<=			16'h0713;
		end
		32'h0000518E: begin
				q			<=			16'h05B6;
		end
		32'h00005190: begin
				q			<=			16'hF06F;
		end
		32'h00005192: begin
				q			<=			16'hFADF;
		end
		32'h00005194: begin
				q			<=			16'h0713;
		end
		32'h00005196: begin
				q			<=			16'h0540;
		end
		32'h00005198: begin
				q			<=			16'h6863;
		end
		32'h0000519A: begin
				q			<=			16'h00C7;
		end
		32'h0000519C: begin
				q			<=			16'hD713;
		end
		32'h0000519E: begin
				q			<=			16'h00C7;
		end
		32'h000051A0: begin
				q			<=			16'h0713;
		end
		32'h000051A2: begin
				q			<=			16'h06E7;
		end
		32'h000051A4: begin
				q			<=			16'hF06F;
		end
		32'h000051A6: begin
				q			<=			16'hF99F;
		end
		32'h000051A8: begin
				q			<=			16'h0713;
		end
		32'h000051AA: begin
				q			<=			16'h1540;
		end
		32'h000051AC: begin
				q			<=			16'h6863;
		end
		32'h000051AE: begin
				q			<=			16'h00C7;
		end
		32'h000051B0: begin
				q			<=			16'hD713;
		end
		32'h000051B2: begin
				q			<=			16'h00F7;
		end
		32'h000051B4: begin
				q			<=			16'h0713;
		end
		32'h000051B6: begin
				q			<=			16'h0777;
		end
		32'h000051B8: begin
				q			<=			16'hF06F;
		end
		32'h000051BA: begin
				q			<=			16'hF85F;
		end
		32'h000051BC: begin
				q			<=			16'h0593;
		end
		32'h000051BE: begin
				q			<=			16'h5540;
		end
		32'h000051C0: begin
				q			<=			16'h0713;
		end
		32'h000051C2: begin
				q			<=			16'h07E0;
		end
		32'h000051C4: begin
				q			<=			16'hECE3;
		end
		32'h000051C6: begin
				q			<=			16'hF6C5;
		end
		32'h000051C8: begin
				q			<=			16'hD713;
		end
		32'h000051CA: begin
				q			<=			16'h0127;
		end
		32'h000051CC: begin
				q			<=			16'h0713;
		end
		32'h000051CE: begin
				q			<=			16'h07C7;
		end
		32'h000051D0: begin
				q			<=			16'hF06F;
		end
		32'h000051D2: begin
				q			<=			16'hF6DF;
		end
		32'h000051D4: begin
				q			<=			16'h2603;
		end
		32'h000051D6: begin
				q			<=			16'h0086;
		end
		32'h000051D8: begin
				q			<=			16'h8863;
		end
		32'h000051DA: begin
				q			<=			16'h00C5;
		end
		32'h000051DC: begin
				q			<=			16'h2703;
		end
		32'h000051DE: begin
				q			<=			16'h0046;
		end
		32'h000051E0: begin
				q			<=			16'h7713;
		end
		32'h000051E2: begin
				q			<=			16'hFFC7;
		end
		32'h000051E4: begin
				q			<=			16'hE8E3;
		end
		32'h000051E6: begin
				q			<=			16'hFEE7;
		end
		32'h000051E8: begin
				q			<=			16'h2583;
		end
		32'h000051EA: begin
				q			<=			16'h00C6;
		end
		32'h000051EC: begin
				q			<=			16'hF06F;
		end
		32'h000051EE: begin
				q			<=			16'hF85F;
		end
		32'h000051F0: begin
				q			<=			16'h8067;
		end
		32'h000051F2: begin
				q			<=			16'h0000;
		end
		32'h000051F4: begin
				q			<=			16'h0000;
		end
		32'h000051F6: begin
				q			<=			16'h0000;
		end
		32'h000051F8: begin
				q			<=			16'h0793;
		end
		32'h000051FA: begin
				q			<=			16'h0145;
		end
		32'h000051FC: begin
				q			<=			16'h0513;
		end
		32'h000051FE: begin
				q			<=			16'h0025;
		end
		32'h00005200: begin
				q			<=			16'h1F23;
		end
		32'h00005202: begin
				q			<=			16'hFE05;
		end
		32'h00005204: begin
				q			<=			16'h1CE3;
		end
		32'h00005206: begin
				q			<=			16'hFEF5;
		end
		32'h00005208: begin
				q			<=			16'h8067;
		end
		32'h0000520A: begin
				q			<=			16'h0000;
		end
		32'h0000520C: begin
				q			<=			16'h0793;
		end
		32'h0000520E: begin
				q			<=			16'h0145;
		end
		32'h00005210: begin
				q			<=			16'h0513;
		end
		32'h00005212: begin
				q			<=			16'h0025;
		end
		32'h00005214: begin
				q			<=			16'h5703;
		end
		32'h00005216: begin
				q			<=			16'hFFE5;
		end
		32'h00005218: begin
				q			<=			16'h8593;
		end
		32'h0000521A: begin
				q			<=			16'h0025;
		end
		32'h0000521C: begin
				q			<=			16'h9F23;
		end
		32'h0000521E: begin
				q			<=			16'hFEE5;
		end
		32'h00005220: begin
				q			<=			16'h98E3;
		end
		32'h00005222: begin
				q			<=			16'hFEA7;
		end
		32'h00005224: begin
				q			<=			16'h8067;
		end
		32'h00005226: begin
				q			<=			16'h0000;
		end
		32'h00005228: begin
				q			<=			16'h0793;
		end
		32'h0000522A: begin
				q			<=			16'h01A5;
		end
		32'h0000522C: begin
				q			<=			16'h0513;
		end
		32'h0000522E: begin
				q			<=			16'h0025;
		end
		32'h00005230: begin
				q			<=			16'h1F23;
		end
		32'h00005232: begin
				q			<=			16'hFE05;
		end
		32'h00005234: begin
				q			<=			16'h1CE3;
		end
		32'h00005236: begin
				q			<=			16'hFEF5;
		end
		32'h00005238: begin
				q			<=			16'h8067;
		end
		32'h0000523A: begin
				q			<=			16'h0000;
		end
		32'h0000523C: begin
				q			<=			16'h0713;
		end
		32'h0000523E: begin
				q			<=			16'h0185;
		end
		32'h00005240: begin
				q			<=			16'h8793;
		end
		32'h00005242: begin
				q			<=			16'h0005;
		end
		32'h00005244: begin
				q			<=			16'h0513;
		end
		32'h00005246: begin
				q			<=			16'h0025;
		end
		32'h00005248: begin
				q			<=			16'h5683;
		end
		32'h0000524A: begin
				q			<=			16'hFFE5;
		end
		32'h0000524C: begin
				q			<=			16'h8793;
		end
		32'h0000524E: begin
				q			<=			16'h0027;
		end
		32'h00005250: begin
				q			<=			16'h9F23;
		end
		32'h00005252: begin
				q			<=			16'hFED7;
		end
		32'h00005254: begin
				q			<=			16'h18E3;
		end
		32'h00005256: begin
				q			<=			16'hFEA7;
		end
		32'h00005258: begin
				q			<=			16'h9C23;
		end
		32'h0000525A: begin
				q			<=			16'h0005;
		end
		32'h0000525C: begin
				q			<=			16'h8067;
		end
		32'h0000525E: begin
				q			<=			16'h0000;
		end
		32'h00005260: begin
				q			<=			16'h0793;
		end
		32'h00005262: begin
				q			<=			16'h0045;
		end
		32'h00005264: begin
				q			<=			16'h8593;
		end
		32'h00005266: begin
				q			<=			16'h0045;
		end
		32'h00005268: begin
				q			<=			16'h0513;
		end
		32'h0000526A: begin
				q			<=			16'h01A5;
		end
		32'h0000526C: begin
				q			<=			16'h8793;
		end
		32'h0000526E: begin
				q			<=			16'h0027;
		end
		32'h00005270: begin
				q			<=			16'h8593;
		end
		32'h00005272: begin
				q			<=			16'h0025;
		end
		32'h00005274: begin
				q			<=			16'hD683;
		end
		32'h00005276: begin
				q			<=			16'hFFE7;
		end
		32'h00005278: begin
				q			<=			16'hD703;
		end
		32'h0000527A: begin
				q			<=			16'hFFE5;
		end
		32'h0000527C: begin
				q			<=			16'h9863;
		end
		32'h0000527E: begin
				q			<=			16'h00E6;
		end
		32'h00005280: begin
				q			<=			16'h16E3;
		end
		32'h00005282: begin
				q			<=			16'hFEF5;
		end
		32'h00005284: begin
				q			<=			16'h0513;
		end
		32'h00005286: begin
				q			<=			16'h0000;
		end
		32'h00005288: begin
				q			<=			16'h8067;
		end
		32'h0000528A: begin
				q			<=			16'h0000;
		end
		32'h0000528C: begin
				q			<=			16'h0513;
		end
		32'h0000528E: begin
				q			<=			16'h0010;
		end
		32'h00005290: begin
				q			<=			16'h6463;
		end
		32'h00005292: begin
				q			<=			16'h00D7;
		end
		32'h00005294: begin
				q			<=			16'h0513;
		end
		32'h00005296: begin
				q			<=			16'hFFF0;
		end
		32'h00005298: begin
				q			<=			16'h8067;
		end
		32'h0000529A: begin
				q			<=			16'h0000;
		end
		32'h0000529C: begin
				q			<=			16'h0693;
		end
		32'h0000529E: begin
				q			<=			16'h0045;
		end
		32'h000052A0: begin
				q			<=			16'h0793;
		end
		32'h000052A2: begin
				q			<=			16'h0000;
		end
		32'h000052A4: begin
				q			<=			16'h0513;
		end
		32'h000052A6: begin
				q			<=			16'h01A5;
		end
		32'h000052A8: begin
				q			<=			16'h8637;
		end
		32'h000052AA: begin
				q			<=			16'hFFFF;
		end
		32'h000052AC: begin
				q			<=			16'hD703;
		end
		32'h000052AE: begin
				q			<=			16'h0006;
		end
		32'h000052B0: begin
				q			<=			16'h7593;
		end
		32'h000052B2: begin
				q			<=			16'h0017;
		end
		32'h000052B4: begin
				q			<=			16'h8463;
		end
		32'h000052B6: begin
				q			<=			16'h0005;
		end
		32'h000052B8: begin
				q			<=			16'hE793;
		end
		32'h000052BA: begin
				q			<=			16'h0017;
		end
		32'h000052BC: begin
				q			<=			16'hF593;
		end
		32'h000052BE: begin
				q			<=			16'h0027;
		end
		32'h000052C0: begin
				q			<=			16'h5713;
		end
		32'h000052C2: begin
				q			<=			16'h0017;
		end
		32'h000052C4: begin
				q			<=			16'h9063;
		end
		32'h000052C6: begin
				q			<=			16'h0205;
		end
		32'h000052C8: begin
				q			<=			16'h9793;
		end
		32'h000052CA: begin
				q			<=			16'h0017;
		end
		32'h000052CC: begin
				q			<=			16'h9023;
		end
		32'h000052CE: begin
				q			<=			16'h00E6;
		end
		32'h000052D0: begin
				q			<=			16'h9793;
		end
		32'h000052D2: begin
				q			<=			16'h0107;
		end
		32'h000052D4: begin
				q			<=			16'h8693;
		end
		32'h000052D6: begin
				q			<=			16'h0026;
		end
		32'h000052D8: begin
				q			<=			16'hD793;
		end
		32'h000052DA: begin
				q			<=			16'h0107;
		end
		32'h000052DC: begin
				q			<=			16'h18E3;
		end
		32'h000052DE: begin
				q			<=			16'hFCD5;
		end
		32'h000052E0: begin
				q			<=			16'h8067;
		end
		32'h000052E2: begin
				q			<=			16'h0000;
		end
		32'h000052E4: begin
				q			<=			16'h6733;
		end
		32'h000052E6: begin
				q			<=			16'h00C7;
		end
		32'h000052E8: begin
				q			<=			16'hF06F;
		end
		32'h000052EA: begin
				q			<=			16'hFE1F;
		end
		32'h000052EC: begin
				q			<=			16'h0693;
		end
		32'h000052EE: begin
				q			<=			16'h0165;
		end
		32'h000052F0: begin
				q			<=			16'h0713;
		end
		32'h000052F2: begin
				q			<=			16'h0000;
		end
		32'h000052F4: begin
				q			<=			16'hD783;
		end
		32'h000052F6: begin
				q			<=			16'h0026;
		end
		32'h000052F8: begin
				q			<=			16'h9613;
		end
		32'h000052FA: begin
				q			<=			16'h0107;
		end
		32'h000052FC: begin
				q			<=			16'h5613;
		end
		32'h000052FE: begin
				q			<=			16'h4106;
		end
		32'h00005300: begin
				q			<=			16'h5463;
		end
		32'h00005302: begin
				q			<=			16'h0006;
		end
		32'h00005304: begin
				q			<=			16'h6713;
		end
		32'h00005306: begin
				q			<=			16'h0017;
		end
		32'h00005308: begin
				q			<=			16'h9793;
		end
		32'h0000530A: begin
				q			<=			16'h0017;
		end
		32'h0000530C: begin
				q			<=			16'h9793;
		end
		32'h0000530E: begin
				q			<=			16'h0107;
		end
		32'h00005310: begin
				q			<=			16'h7613;
		end
		32'h00005312: begin
				q			<=			16'h0027;
		end
		32'h00005314: begin
				q			<=			16'hD793;
		end
		32'h00005316: begin
				q			<=			16'h0107;
		end
		32'h00005318: begin
				q			<=			16'h1063;
		end
		32'h0000531A: begin
				q			<=			16'h0206;
		end
		32'h0000531C: begin
				q			<=			16'h1713;
		end
		32'h0000531E: begin
				q			<=			16'h0017;
		end
		32'h00005320: begin
				q			<=			16'h9123;
		end
		32'h00005322: begin
				q			<=			16'h00F6;
		end
		32'h00005324: begin
				q			<=			16'h1713;
		end
		32'h00005326: begin
				q			<=			16'h0107;
		end
		32'h00005328: begin
				q			<=			16'h8693;
		end
		32'h0000532A: begin
				q			<=			16'hFFE6;
		end
		32'h0000532C: begin
				q			<=			16'h5713;
		end
		32'h0000532E: begin
				q			<=			16'h0107;
		end
		32'h00005330: begin
				q			<=			16'h12E3;
		end
		32'h00005332: begin
				q			<=			16'hFCD5;
		end
		32'h00005334: begin
				q			<=			16'h8067;
		end
		32'h00005336: begin
				q			<=			16'h0000;
		end
		32'h00005338: begin
				q			<=			16'hE793;
		end
		32'h0000533A: begin
				q			<=			16'h0017;
		end
		32'h0000533C: begin
				q			<=			16'hF06F;
		end
		32'h0000533E: begin
				q			<=			16'hFE1F;
		end
		32'h00005340: begin
				q			<=			16'h0793;
		end
		32'h00005342: begin
				q			<=			16'h0045;
		end
		32'h00005344: begin
				q			<=			16'h0713;
		end
		32'h00005346: begin
				q			<=			16'h0000;
		end
		32'h00005348: begin
				q			<=			16'h0513;
		end
		32'h0000534A: begin
				q			<=			16'h01A5;
		end
		32'h0000534C: begin
				q			<=			16'hD683;
		end
		32'h0000534E: begin
				q			<=			16'h0007;
		end
		32'h00005350: begin
				q			<=			16'h8793;
		end
		32'h00005352: begin
				q			<=			16'h0027;
		end
		32'h00005354: begin
				q			<=			16'hD613;
		end
		32'h00005356: begin
				q			<=			16'h0086;
		end
		32'h00005358: begin
				q			<=			16'h6733;
		end
		32'h0000535A: begin
				q			<=			16'h00C7;
		end
		32'h0000535C: begin
				q			<=			16'h9F23;
		end
		32'h0000535E: begin
				q			<=			16'hFEE7;
		end
		32'h00005360: begin
				q			<=			16'h9713;
		end
		32'h00005362: begin
				q			<=			16'h0086;
		end
		32'h00005364: begin
				q			<=			16'h1713;
		end
		32'h00005366: begin
				q			<=			16'h0107;
		end
		32'h00005368: begin
				q			<=			16'h5713;
		end
		32'h0000536A: begin
				q			<=			16'h0107;
		end
		32'h0000536C: begin
				q			<=			16'h10E3;
		end
		32'h0000536E: begin
				q			<=			16'hFEF5;
		end
		32'h00005370: begin
				q			<=			16'h8067;
		end
		32'h00005372: begin
				q			<=			16'h0000;
		end
		32'h00005374: begin
				q			<=			16'h0793;
		end
		32'h00005376: begin
				q			<=			16'h0165;
		end
		32'h00005378: begin
				q			<=			16'h0713;
		end
		32'h0000537A: begin
				q			<=			16'h0000;
		end
		32'h0000537C: begin
				q			<=			16'hD683;
		end
		32'h0000537E: begin
				q			<=			16'h0027;
		end
		32'h00005380: begin
				q			<=			16'h8793;
		end
		32'h00005382: begin
				q			<=			16'hFFE7;
		end
		32'h00005384: begin
				q			<=			16'h9613;
		end
		32'h00005386: begin
				q			<=			16'h0086;
		end
		32'h00005388: begin
				q			<=			16'h6733;
		end
		32'h0000538A: begin
				q			<=			16'h00C7;
		end
		32'h0000538C: begin
				q			<=			16'h9223;
		end
		32'h0000538E: begin
				q			<=			16'h00E7;
		end
		32'h00005390: begin
				q			<=			16'hD713;
		end
		32'h00005392: begin
				q			<=			16'h0086;
		end
		32'h00005394: begin
				q			<=			16'h14E3;
		end
		32'h00005396: begin
				q			<=			16'hFEF5;
		end
		32'h00005398: begin
				q			<=			16'h8067;
		end
		32'h0000539A: begin
				q			<=			16'h0000;
		end
		32'h0000539C: begin
				q			<=			16'h0793;
		end
		32'h0000539E: begin
				q			<=			16'h0045;
		end
		32'h000053A0: begin
				q			<=			16'h0713;
		end
		32'h000053A2: begin
				q			<=			16'h0185;
		end
		32'h000053A4: begin
				q			<=			16'h8793;
		end
		32'h000053A6: begin
				q			<=			16'h0027;
		end
		32'h000053A8: begin
				q			<=			16'hD683;
		end
		32'h000053AA: begin
				q			<=			16'h0007;
		end
		32'h000053AC: begin
				q			<=			16'h9F23;
		end
		32'h000053AE: begin
				q			<=			16'hFED7;
		end
		32'h000053B0: begin
				q			<=			16'h1AE3;
		end
		32'h000053B2: begin
				q			<=			16'hFEF7;
		end
		32'h000053B4: begin
				q			<=			16'h1C23;
		end
		32'h000053B6: begin
				q			<=			16'h0005;
		end
		32'h000053B8: begin
				q			<=			16'h8067;
		end
		32'h000053BA: begin
				q			<=			16'h0000;
		end
		32'h000053BC: begin
				q			<=			16'h0793;
		end
		32'h000053BE: begin
				q			<=			16'h0185;
		end
		32'h000053C0: begin
				q			<=			16'h0713;
		end
		32'h000053C2: begin
				q			<=			16'h01A5;
		end
		32'h000053C4: begin
				q			<=			16'h0693;
		end
		32'h000053C6: begin
				q			<=			16'h0045;
		end
		32'h000053C8: begin
				q			<=			16'h8793;
		end
		32'h000053CA: begin
				q			<=			16'hFFE7;
		end
		32'h000053CC: begin
				q			<=			16'hD603;
		end
		32'h000053CE: begin
				q			<=			16'h0007;
		end
		32'h000053D0: begin
				q			<=			16'h0713;
		end
		32'h000053D2: begin
				q			<=			16'hFFE7;
		end
		32'h000053D4: begin
				q			<=			16'h1023;
		end
		32'h000053D6: begin
				q			<=			16'h00C7;
		end
		32'h000053D8: begin
				q			<=			16'h98E3;
		end
		32'h000053DA: begin
				q			<=			16'hFEF6;
		end
		32'h000053DC: begin
				q			<=			16'h1223;
		end
		32'h000053DE: begin
				q			<=			16'h0005;
		end
		32'h000053E0: begin
				q			<=			16'h8067;
		end
		32'h000053E2: begin
				q			<=			16'h0000;
		end
		32'h000053E4: begin
				q			<=			16'h8593;
		end
		32'h000053E6: begin
				q			<=			16'h0185;
		end
		32'h000053E8: begin
				q			<=			16'h0713;
		end
		32'h000053EA: begin
				q			<=			16'h0165;
		end
		32'h000053EC: begin
				q			<=			16'h0693;
		end
		32'h000053EE: begin
				q			<=			16'h0000;
		end
		32'h000053F0: begin
				q			<=			16'h5783;
		end
		32'h000053F2: begin
				q			<=			16'h0027;
		end
		32'h000053F4: begin
				q			<=			16'hD603;
		end
		32'h000053F6: begin
				q			<=			16'h0005;
		end
		32'h000053F8: begin
				q			<=			16'h0713;
		end
		32'h000053FA: begin
				q			<=			16'hFFE7;
		end
		32'h000053FC: begin
				q			<=			16'h8593;
		end
		32'h000053FE: begin
				q			<=			16'hFFE5;
		end
		32'h00005400: begin
				q			<=			16'h87B3;
		end
		32'h00005402: begin
				q			<=			16'h00C7;
		end
		32'h00005404: begin
				q			<=			16'h87B3;
		end
		32'h00005406: begin
				q			<=			16'h00D7;
		end
		32'h00005408: begin
				q			<=			16'h9123;
		end
		32'h0000540A: begin
				q			<=			16'h00F5;
		end
		32'h0000540C: begin
				q			<=			16'hD793;
		end
		32'h0000540E: begin
				q			<=			16'h0107;
		end
		32'h00005410: begin
				q			<=			16'hF693;
		end
		32'h00005412: begin
				q			<=			16'h0017;
		end
		32'h00005414: begin
				q			<=			16'h1EE3;
		end
		32'h00005416: begin
				q			<=			16'hFCE5;
		end
		32'h00005418: begin
				q			<=			16'h8067;
		end
		32'h0000541A: begin
				q			<=			16'h0000;
		end
		32'h0000541C: begin
				q			<=			16'h8593;
		end
		32'h0000541E: begin
				q			<=			16'h0185;
		end
		32'h00005420: begin
				q			<=			16'h0713;
		end
		32'h00005422: begin
				q			<=			16'h0165;
		end
		32'h00005424: begin
				q			<=			16'h0693;
		end
		32'h00005426: begin
				q			<=			16'h0000;
		end
		32'h00005428: begin
				q			<=			16'hD783;
		end
		32'h0000542A: begin
				q			<=			16'h0005;
		end
		32'h0000542C: begin
				q			<=			16'h5603;
		end
		32'h0000542E: begin
				q			<=			16'h0027;
		end
		32'h00005430: begin
				q			<=			16'h0713;
		end
		32'h00005432: begin
				q			<=			16'hFFE7;
		end
		32'h00005434: begin
				q			<=			16'h8593;
		end
		32'h00005436: begin
				q			<=			16'hFFE5;
		end
		32'h00005438: begin
				q			<=			16'h87B3;
		end
		32'h0000543A: begin
				q			<=			16'h40C7;
		end
		32'h0000543C: begin
				q			<=			16'h87B3;
		end
		32'h0000543E: begin
				q			<=			16'h40D7;
		end
		32'h00005440: begin
				q			<=			16'h9123;
		end
		32'h00005442: begin
				q			<=			16'h00F5;
		end
		32'h00005444: begin
				q			<=			16'hD793;
		end
		32'h00005446: begin
				q			<=			16'h0107;
		end
		32'h00005448: begin
				q			<=			16'hF693;
		end
		32'h0000544A: begin
				q			<=			16'h0017;
		end
		32'h0000544C: begin
				q			<=			16'h1EE3;
		end
		32'h0000544E: begin
				q			<=			16'hFCE5;
		end
		32'h00005450: begin
				q			<=			16'h8067;
		end
		32'h00005452: begin
				q			<=			16'h0000;
		end
		32'h00005454: begin
				q			<=			16'h0113;
		end
		32'h00005456: begin
				q			<=			16'hFE01;
		end
		32'h00005458: begin
				q			<=			16'h0337;
		end
		32'h0000545A: begin
				q			<=			16'h0001;
		end
		32'h0000545C: begin
				q			<=			16'h8893;
		end
		32'h0000545E: begin
				q			<=			16'h0185;
		end
		32'h00005460: begin
				q			<=			16'h1D23;
		end
		32'h00005462: begin
				q			<=			16'h0001;
		end
		32'h00005464: begin
				q			<=			16'h1E23;
		end
		32'h00005466: begin
				q			<=			16'h0001;
		end
		32'h00005468: begin
				q			<=			16'h8593;
		end
		32'h0000546A: begin
				q			<=			16'h0045;
		end
		32'h0000546C: begin
				q			<=			16'h0693;
		end
		32'h0000546E: begin
				q			<=			16'h01C1;
		end
		32'h00005470: begin
				q			<=			16'h0313;
		end
		32'h00005472: begin
				q			<=			16'hFFF3;
		end
		32'h00005474: begin
				q			<=			16'hD703;
		end
		32'h00005476: begin
				q			<=			16'h0008;
		end
		32'h00005478: begin
				q			<=			16'h8693;
		end
		32'h0000547A: begin
				q			<=			16'hFFE6;
		end
		32'h0000547C: begin
				q			<=			16'h8893;
		end
		32'h0000547E: begin
				q			<=			16'hFFE8;
		end
		32'h00005480: begin
				q			<=			16'h1C63;
		end
		32'h00005482: begin
				q			<=			16'h0207;
		end
		32'h00005484: begin
				q			<=			16'h9F23;
		end
		32'h00005486: begin
				q			<=			16'hFE06;
		end
		32'h00005488: begin
				q			<=			16'h96E3;
		end
		32'h0000548A: begin
				q			<=			16'hFF15;
		end
		32'h0000548C: begin
				q			<=			16'h0793;
		end
		32'h0000548E: begin
				q			<=			16'h0040;
		end
		32'h00005490: begin
				q			<=			16'h0713;
		end
		32'h00005492: begin
				q			<=			16'h01A0;
		end
		32'h00005494: begin
				q			<=			16'h0593;
		end
		32'h00005496: begin
				q			<=			16'h0041;
		end
		32'h00005498: begin
				q			<=			16'h85B3;
		end
		32'h0000549A: begin
				q			<=			16'h00F5;
		end
		32'h0000549C: begin
				q			<=			16'hD583;
		end
		32'h0000549E: begin
				q			<=			16'h0005;
		end
		32'h000054A0: begin
				q			<=			16'h06B3;
		end
		32'h000054A2: begin
				q			<=			16'h00F6;
		end
		32'h000054A4: begin
				q			<=			16'h8793;
		end
		32'h000054A6: begin
				q			<=			16'h0027;
		end
		32'h000054A8: begin
				q			<=			16'h9023;
		end
		32'h000054AA: begin
				q			<=			16'h00B6;
		end
		32'h000054AC: begin
				q			<=			16'h94E3;
		end
		32'h000054AE: begin
				q			<=			16'hFEE7;
		end
		32'h000054B0: begin
				q			<=			16'h0113;
		end
		32'h000054B2: begin
				q			<=			16'h0201;
		end
		32'h000054B4: begin
				q			<=			16'h8067;
		end
		32'h000054B6: begin
				q			<=			16'h0000;
		end
		32'h000054B8: begin
				q			<=			16'h0733;
		end
		32'h000054BA: begin
				q			<=			16'h02A7;
		end
		32'h000054BC: begin
				q			<=			16'hD803;
		end
		32'h000054BE: begin
				q			<=			16'h0026;
		end
		32'h000054C0: begin
				q			<=			16'h77B3;
		end
		32'h000054C2: begin
				q			<=			16'h0067;
		end
		32'h000054C4: begin
				q			<=			16'h87B3;
		end
		32'h000054C6: begin
				q			<=			16'h0107;
		end
		32'h000054C8: begin
				q			<=			16'hD813;
		end
		32'h000054CA: begin
				q			<=			16'h0107;
		end
		32'h000054CC: begin
				q			<=			16'h9123;
		end
		32'h000054CE: begin
				q			<=			16'h00F6;
		end
		32'h000054D0: begin
				q			<=			16'h5793;
		end
		32'h000054D2: begin
				q			<=			16'h0107;
		end
		32'h000054D4: begin
				q			<=			16'hD703;
		end
		32'h000054D6: begin
				q			<=			16'h0006;
		end
		32'h000054D8: begin
				q			<=			16'h87B3;
		end
		32'h000054DA: begin
				q			<=			16'h00E7;
		end
		32'h000054DC: begin
				q			<=			16'h87B3;
		end
		32'h000054DE: begin
				q			<=			16'h0107;
		end
		32'h000054E0: begin
				q			<=			16'h9023;
		end
		32'h000054E2: begin
				q			<=			16'h00F6;
		end
		32'h000054E4: begin
				q			<=			16'hD793;
		end
		32'h000054E6: begin
				q			<=			16'h0107;
		end
		32'h000054E8: begin
				q			<=			16'h9F23;
		end
		32'h000054EA: begin
				q			<=			16'hFEF6;
		end
		32'h000054EC: begin
				q			<=			16'hF06F;
		end
		32'h000054EE: begin
				q			<=			16'hF9DF;
		end
		32'h000054F0: begin
				q			<=			16'h5783;
		end
		32'h000054F2: begin
				q			<=			16'h0125;
		end
		32'h000054F4: begin
				q			<=			16'hC793;
		end
		32'h000054F6: begin
				q			<=			16'hFFF7;
		end
		32'h000054F8: begin
				q			<=			16'h9713;
		end
		32'h000054FA: begin
				q			<=			16'h0117;
		end
		32'h000054FC: begin
				q			<=			16'h1C63;
		end
		32'h000054FE: begin
				q			<=			16'h0007;
		end
		32'h00005500: begin
				q			<=			16'h0793;
		end
		32'h00005502: begin
				q			<=			16'h0125;
		end
		32'h00005504: begin
				q			<=			16'h0513;
		end
		32'h00005506: begin
				q			<=			16'h0025;
		end
		32'h00005508: begin
				q			<=			16'h5703;
		end
		32'h0000550A: begin
				q			<=			16'hFFE5;
		end
		32'h0000550C: begin
				q			<=			16'h1863;
		end
		32'h0000550E: begin
				q			<=			16'h0007;
		end
		32'h00005510: begin
				q			<=			16'h9AE3;
		end
		32'h00005512: begin
				q			<=			16'hFEA7;
		end
		32'h00005514: begin
				q			<=			16'h0513;
		end
		32'h00005516: begin
				q			<=			16'h0000;
		end
		32'h00005518: begin
				q			<=			16'h8067;
		end
		32'h0000551A: begin
				q			<=			16'h0000;
		end
		32'h0000551C: begin
				q			<=			16'h0513;
		end
		32'h0000551E: begin
				q			<=			16'h0010;
		end
		32'h00005520: begin
				q			<=			16'h8067;
		end
		32'h00005522: begin
				q			<=			16'h0000;
		end
		32'h00005524: begin
				q			<=			16'h0113;
		end
		32'h00005526: begin
				q			<=			16'hFF01;
		end
		32'h00005528: begin
				q			<=			16'h2423;
		end
		32'h0000552A: begin
				q			<=			16'h0081;
		end
		32'h0000552C: begin
				q			<=			16'h2623;
		end
		32'h0000552E: begin
				q			<=			16'h0011;
		end
		32'h00005530: begin
				q			<=			16'h0413;
		end
		32'h00005532: begin
				q			<=			16'h0005;
		end
		32'h00005534: begin
				q			<=			16'h0097;
		end
		32'h00005536: begin
				q			<=			16'h0000;
		end
		32'h00005538: begin
				q			<=			16'h80E7;
		end
		32'h0000553A: begin
				q			<=			16'hFBC0;
		end
		32'h0000553C: begin
				q			<=			16'h1E63;
		end
		32'h0000553E: begin
				q			<=			16'h0005;
		end
		32'h00005540: begin
				q			<=			16'h1503;
		end
		32'h00005542: begin
				q			<=			16'h0124;
		end
		32'h00005544: begin
				q			<=			16'h5513;
		end
		32'h00005546: begin
				q			<=			16'h01F5;
		end
		32'h00005548: begin
				q			<=			16'h2083;
		end
		32'h0000554A: begin
				q			<=			16'h00C1;
		end
		32'h0000554C: begin
				q			<=			16'h2403;
		end
		32'h0000554E: begin
				q			<=			16'h0081;
		end
		32'h00005550: begin
				q			<=			16'h0113;
		end
		32'h00005552: begin
				q			<=			16'h0101;
		end
		32'h00005554: begin
				q			<=			16'h8067;
		end
		32'h00005556: begin
				q			<=			16'h0000;
		end
		32'h00005558: begin
				q			<=			16'h0513;
		end
		32'h0000555A: begin
				q			<=			16'h0000;
		end
		32'h0000555C: begin
				q			<=			16'hF06F;
		end
		32'h0000555E: begin
				q			<=			16'hFEDF;
		end
		32'h00005560: begin
				q			<=			16'h1783;
		end
		32'h00005562: begin
				q			<=			16'h0125;
		end
		32'h00005564: begin
				q			<=			16'h0113;
		end
		32'h00005566: begin
				q			<=			16'hFF01;
		end
		32'h00005568: begin
				q			<=			16'h2623;
		end
		32'h0000556A: begin
				q			<=			16'h0011;
		end
		32'h0000556C: begin
				q			<=			16'h2423;
		end
		32'h0000556E: begin
				q			<=			16'h0081;
		end
		32'h00005570: begin
				q			<=			16'h2223;
		end
		32'h00005572: begin
				q			<=			16'h0091;
		end
		32'h00005574: begin
				q			<=			16'h2023;
		end
		32'h00005576: begin
				q			<=			16'h0121;
		end
		32'h00005578: begin
				q			<=			16'hD863;
		end
		32'h0000557A: begin
				q			<=			16'h0607;
		end
		32'h0000557C: begin
				q			<=			16'h0793;
		end
		32'h0000557E: begin
				q			<=			16'hFFF0;
		end
		32'h00005580: begin
				q			<=			16'h9023;
		end
		32'h00005582: begin
				q			<=			16'h00F5;
		end
		32'h00005584: begin
				q			<=			16'h5703;
		end
		32'h00005586: begin
				q			<=			16'h0125;
		end
		32'h00005588: begin
				q			<=			16'h87B7;
		end
		32'h0000558A: begin
				q			<=			16'h0000;
		end
		32'h0000558C: begin
				q			<=			16'h8793;
		end
		32'h0000558E: begin
				q			<=			16'hFFF7;
		end
		32'h00005590: begin
				q			<=			16'hF733;
		end
		32'h00005592: begin
				q			<=			16'h00E7;
		end
		32'h00005594: begin
				q			<=			16'h9123;
		end
		32'h00005596: begin
				q			<=			16'h00E5;
		end
		32'h00005598: begin
				q			<=			16'h0913;
		end
		32'h0000559A: begin
				q			<=			16'h0105;
		end
		32'h0000559C: begin
				q			<=			16'h1663;
		end
		32'h0000559E: begin
				q			<=			16'h06F7;
		end
		32'h000055A0: begin
				q			<=			16'h8413;
		end
		32'h000055A2: begin
				q			<=			16'h0005;
		end
		32'h000055A4: begin
				q			<=			16'h0493;
		end
		32'h000055A6: begin
				q			<=			16'h0005;
		end
		32'h000055A8: begin
				q			<=			16'hF0EF;
		end
		32'h000055AA: begin
				q			<=			16'hF49F;
		end
		32'h000055AC: begin
				q			<=			16'h0263;
		end
		32'h000055AE: begin
				q			<=			16'h0405;
		end
		32'h000055B0: begin
				q			<=			16'h0793;
		end
		32'h000055B2: begin
				q			<=			16'h0064;
		end
		32'h000055B4: begin
				q			<=			16'h1223;
		end
		32'h000055B6: begin
				q			<=			16'h0004;
		end
		32'h000055B8: begin
				q			<=			16'h8513;
		end
		32'h000055BA: begin
				q			<=			16'hFFC4;
		end
		32'h000055BC: begin
				q			<=			16'h0913;
		end
		32'h000055BE: begin
				q			<=			16'hFFE9;
		end
		32'h000055C0: begin
				q			<=			16'h5703;
		end
		32'h000055C2: begin
				q			<=			16'h0029;
		end
		32'h000055C4: begin
				q			<=			16'h8793;
		end
		32'h000055C6: begin
				q			<=			16'h0027;
		end
		32'h000055C8: begin
				q			<=			16'h9F23;
		end
		32'h000055CA: begin
				q			<=			16'hFEE7;
		end
		32'h000055CC: begin
				q			<=			16'h18E3;
		end
		32'h000055CE: begin
				q			<=			16'hFEA9;
		end
		32'h000055D0: begin
				q			<=			16'h2083;
		end
		32'h000055D2: begin
				q			<=			16'h00C1;
		end
		32'h000055D4: begin
				q			<=			16'h2403;
		end
		32'h000055D6: begin
				q			<=			16'h0081;
		end
		32'h000055D8: begin
				q			<=			16'h2483;
		end
		32'h000055DA: begin
				q			<=			16'h0041;
		end
		32'h000055DC: begin
				q			<=			16'h2903;
		end
		32'h000055DE: begin
				q			<=			16'h0001;
		end
		32'h000055E0: begin
				q			<=			16'h0113;
		end
		32'h000055E2: begin
				q			<=			16'h0101;
		end
		32'h000055E4: begin
				q			<=			16'h8067;
		end
		32'h000055E6: begin
				q			<=			16'h0000;
		end
		32'h000055E8: begin
				q			<=			16'h9023;
		end
		32'h000055EA: begin
				q			<=			16'h0005;
		end
		32'h000055EC: begin
				q			<=			16'hF06F;
		end
		32'h000055EE: begin
				q			<=			16'hF99F;
		end
		32'h000055F0: begin
				q			<=			16'h0793;
		end
		32'h000055F2: begin
				q			<=			16'h0044;
		end
		32'h000055F4: begin
				q			<=			16'h0593;
		end
		32'h000055F6: begin
				q			<=			16'h01A4;
		end
		32'h000055F8: begin
				q			<=			16'h8793;
		end
		32'h000055FA: begin
				q			<=			16'h0027;
		end
		32'h000055FC: begin
				q			<=			16'h9F23;
		end
		32'h000055FE: begin
				q			<=			16'hFE07;
		end
		32'h00005600: begin
				q			<=			16'h9CE3;
		end
		32'h00005602: begin
				q			<=			16'hFEB7;
		end
		32'h00005604: begin
				q			<=			16'hF06F;
		end
		32'h00005606: begin
				q			<=			16'hFCDF;
		end
		32'h00005608: begin
				q			<=			16'h8793;
		end
		32'h0000560A: begin
				q			<=			16'h0065;
		end
		32'h0000560C: begin
				q			<=			16'h9223;
		end
		32'h0000560E: begin
				q			<=			16'h0005;
		end
		32'h00005610: begin
				q			<=			16'h0513;
		end
		32'h00005612: begin
				q			<=			16'hFFE5;
		end
		32'h00005614: begin
				q			<=			16'h0913;
		end
		32'h00005616: begin
				q			<=			16'hFFE9;
		end
		32'h00005618: begin
				q			<=			16'h5703;
		end
		32'h0000561A: begin
				q			<=			16'h0029;
		end
		32'h0000561C: begin
				q			<=			16'h8793;
		end
		32'h0000561E: begin
				q			<=			16'h0027;
		end
		32'h00005620: begin
				q			<=			16'h9F23;
		end
		32'h00005622: begin
				q			<=			16'hFEE7;
		end
		32'h00005624: begin
				q			<=			16'h18E3;
		end
		32'h00005626: begin
				q			<=			16'hFEA9;
		end
		32'h00005628: begin
				q			<=			16'h9C23;
		end
		32'h0000562A: begin
				q			<=			16'h0005;
		end
		32'h0000562C: begin
				q			<=			16'hF06F;
		end
		32'h0000562E: begin
				q			<=			16'hFA5F;
		end
		32'h00005630: begin
				q			<=			16'h0113;
		end
		32'h00005632: begin
				q			<=			16'hFB01;
		end
		32'h00005634: begin
				q			<=			16'h2223;
		end
		32'h00005636: begin
				q			<=			16'h0491;
		end
		32'h00005638: begin
				q			<=			16'h2023;
		end
		32'h0000563A: begin
				q			<=			16'h0521;
		end
		32'h0000563C: begin
				q			<=			16'h2623;
		end
		32'h0000563E: begin
				q			<=			16'h0411;
		end
		32'h00005640: begin
				q			<=			16'h2423;
		end
		32'h00005642: begin
				q			<=			16'h0481;
		end
		32'h00005644: begin
				q			<=			16'h0913;
		end
		32'h00005646: begin
				q			<=			16'h0005;
		end
		32'h00005648: begin
				q			<=			16'h8493;
		end
		32'h0000564A: begin
				q			<=			16'h0005;
		end
		32'h0000564C: begin
				q			<=			16'h0097;
		end
		32'h0000564E: begin
				q			<=			16'h0000;
		end
		32'h00005650: begin
				q			<=			16'h80E7;
		end
		32'h00005652: begin
				q			<=			16'hEA40;
		end
		32'h00005654: begin
				q			<=			16'h1663;
		end
		32'h00005656: begin
				q			<=			16'h0E05;
		end
		32'h00005658: begin
				q			<=			16'h8513;
		end
		32'h0000565A: begin
				q			<=			16'h0004;
		end
		32'h0000565C: begin
				q			<=			16'h0097;
		end
		32'h0000565E: begin
				q			<=			16'h0000;
		end
		32'h00005660: begin
				q			<=			16'h80E7;
		end
		32'h00005662: begin
				q			<=			16'hE940;
		end
		32'h00005664: begin
				q			<=			16'h0413;
		end
		32'h00005666: begin
				q			<=			16'h0005;
		end
		32'h00005668: begin
				q			<=			16'h1C63;
		end
		32'h0000566A: begin
				q			<=			16'h0C05;
		end
		32'h0000566C: begin
				q			<=			16'h0593;
		end
		32'h0000566E: begin
				q			<=			16'h0081;
		end
		32'h00005670: begin
				q			<=			16'h0513;
		end
		32'h00005672: begin
				q			<=			16'h0009;
		end
		32'h00005674: begin
				q			<=			16'h0097;
		end
		32'h00005676: begin
				q			<=			16'h0000;
		end
		32'h00005678: begin
				q			<=			16'h80E7;
		end
		32'h0000567A: begin
				q			<=			16'hEEC0;
		end
		32'h0000567C: begin
				q			<=			16'h0593;
		end
		32'h0000567E: begin
				q			<=			16'h0241;
		end
		32'h00005680: begin
				q			<=			16'h8513;
		end
		32'h00005682: begin
				q			<=			16'h0004;
		end
		32'h00005684: begin
				q			<=			16'h0097;
		end
		32'h00005686: begin
				q			<=			16'h0000;
		end
		32'h00005688: begin
				q			<=			16'h80E7;
		end
		32'h0000568A: begin
				q			<=			16'hEDC0;
		end
		32'h0000568C: begin
				q			<=			16'h5703;
		end
		32'h0000568E: begin
				q			<=			16'h0081;
		end
		32'h00005690: begin
				q			<=			16'h5783;
		end
		32'h00005692: begin
				q			<=			16'h0241;
		end
		32'h00005694: begin
				q			<=			16'h8063;
		end
		32'h00005696: begin
				q			<=			16'h06E7;
		end
		32'h00005698: begin
				q			<=			16'h0793;
		end
		32'h0000569A: begin
				q			<=			16'h0020;
		end
		32'h0000569C: begin
				q			<=			16'h0693;
		end
		32'h0000569E: begin
				q			<=			16'h0180;
		end
		32'h000056A0: begin
				q			<=			16'h0613;
		end
		32'h000056A2: begin
				q			<=			16'h0081;
		end
		32'h000056A4: begin
				q			<=			16'h0633;
		end
		32'h000056A6: begin
				q			<=			16'h00F6;
		end
		32'h000056A8: begin
				q			<=			16'h5603;
		end
		32'h000056AA: begin
				q			<=			16'h0006;
		end
		32'h000056AC: begin
				q			<=			16'h1C63;
		end
		32'h000056AE: begin
				q			<=			16'h0206;
		end
		32'h000056B0: begin
				q			<=			16'h0613;
		end
		32'h000056B2: begin
				q			<=			16'h0241;
		end
		32'h000056B4: begin
				q			<=			16'h0633;
		end
		32'h000056B6: begin
				q			<=			16'h00F6;
		end
		32'h000056B8: begin
				q			<=			16'h5603;
		end
		32'h000056BA: begin
				q			<=			16'h0006;
		end
		32'h000056BC: begin
				q			<=			16'h1463;
		end
		32'h000056BE: begin
				q			<=			16'h0206;
		end
		32'h000056C0: begin
				q			<=			16'h8793;
		end
		32'h000056C2: begin
				q			<=			16'h0027;
		end
		32'h000056C4: begin
				q			<=			16'h9EE3;
		end
		32'h000056C6: begin
				q			<=			16'hFCD7;
		end
		32'h000056C8: begin
				q			<=			16'h0513;
		end
		32'h000056CA: begin
				q			<=			16'h0004;
		end
		32'h000056CC: begin
				q			<=			16'h2083;
		end
		32'h000056CE: begin
				q			<=			16'h04C1;
		end
		32'h000056D0: begin
				q			<=			16'h2403;
		end
		32'h000056D2: begin
				q			<=			16'h0481;
		end
		32'h000056D4: begin
				q			<=			16'h2483;
		end
		32'h000056D6: begin
				q			<=			16'h0441;
		end
		32'h000056D8: begin
				q			<=			16'h2903;
		end
		32'h000056DA: begin
				q			<=			16'h0401;
		end
		32'h000056DC: begin
				q			<=			16'h0113;
		end
		32'h000056DE: begin
				q			<=			16'h0501;
		end
		32'h000056E0: begin
				q			<=			16'h8067;
		end
		32'h000056E2: begin
				q			<=			16'h0000;
		end
		32'h000056E4: begin
				q			<=			16'h0413;
		end
		32'h000056E6: begin
				q			<=			16'h0010;
		end
		32'h000056E8: begin
				q			<=			16'h00E3;
		end
		32'h000056EA: begin
				q			<=			16'hFE07;
		end
		32'h000056EC: begin
				q			<=			16'h0413;
		end
		32'h000056EE: begin
				q			<=			16'hFFF0;
		end
		32'h000056F0: begin
				q			<=			16'hF06F;
		end
		32'h000056F2: begin
				q			<=			16'hFD9F;
		end
		32'h000056F4: begin
				q			<=			16'h0613;
		end
		32'h000056F6: begin
				q			<=			16'h0010;
		end
		32'h000056F8: begin
				q			<=			16'h8463;
		end
		32'h000056FA: begin
				q			<=			16'h0007;
		end
		32'h000056FC: begin
				q			<=			16'h0613;
		end
		32'h000056FE: begin
				q			<=			16'hFFF0;
		end
		32'h00005700: begin
				q			<=			16'h0793;
		end
		32'h00005702: begin
				q			<=			16'h0000;
		end
		32'h00005704: begin
				q			<=			16'h0593;
		end
		32'h00005706: begin
				q			<=			16'h0180;
		end
		32'h00005708: begin
				q			<=			16'h0713;
		end
		32'h0000570A: begin
				q			<=			16'h0081;
		end
		32'h0000570C: begin
				q			<=			16'h0733;
		end
		32'h0000570E: begin
				q			<=			16'h00F7;
		end
		32'h00005710: begin
				q			<=			16'h5683;
		end
		32'h00005712: begin
				q			<=			16'h0007;
		end
		32'h00005714: begin
				q			<=			16'h0713;
		end
		32'h00005716: begin
				q			<=			16'h0241;
		end
		32'h00005718: begin
				q			<=			16'h0733;
		end
		32'h0000571A: begin
				q			<=			16'h00F7;
		end
		32'h0000571C: begin
				q			<=			16'h5703;
		end
		32'h0000571E: begin
				q			<=			16'h0007;
		end
		32'h00005720: begin
				q			<=			16'h9863;
		end
		32'h00005722: begin
				q			<=			16'h00E6;
		end
		32'h00005724: begin
				q			<=			16'h8793;
		end
		32'h00005726: begin
				q			<=			16'h0027;
		end
		32'h00005728: begin
				q			<=			16'h90E3;
		end
		32'h0000572A: begin
				q			<=			16'hFEB7;
		end
		32'h0000572C: begin
				q			<=			16'hF06F;
		end
		32'h0000572E: begin
				q			<=			16'hF9DF;
		end
		32'h00005730: begin
				q			<=			16'h0413;
		end
		32'h00005732: begin
				q			<=			16'h0006;
		end
		32'h00005734: begin
				q			<=			16'h6AE3;
		end
		32'h00005736: begin
				q			<=			16'hF8D7;
		end
		32'h00005738: begin
				q			<=			16'h0433;
		end
		32'h0000573A: begin
				q			<=			16'h40C0;
		end
		32'h0000573C: begin
				q			<=			16'hF06F;
		end
		32'h0000573E: begin
				q			<=			16'hF8DF;
		end
		32'h00005740: begin
				q			<=			16'h0413;
		end
		32'h00005742: begin
				q			<=			16'hFFE0;
		end
		32'h00005744: begin
				q			<=			16'hF06F;
		end
		32'h00005746: begin
				q			<=			16'hF85F;
		end
		32'h00005748: begin
				q			<=			16'h5783;
		end
		32'h0000574A: begin
				q			<=			16'h0125;
		end
		32'h0000574C: begin
				q			<=			16'hC793;
		end
		32'h0000574E: begin
				q			<=			16'hFFF7;
		end
		32'h00005750: begin
				q			<=			16'h9713;
		end
		32'h00005752: begin
				q			<=			16'h0117;
		end
		32'h00005754: begin
				q			<=			16'h1063;
		end
		32'h00005756: begin
				q			<=			16'h0207;
		end
		32'h00005758: begin
				q			<=			16'h0113;
		end
		32'h0000575A: begin
				q			<=			16'hFF01;
		end
		32'h0000575C: begin
				q			<=			16'h2623;
		end
		32'h0000575E: begin
				q			<=			16'h0011;
		end
		32'h00005760: begin
				q			<=			16'hF0EF;
		end
		32'h00005762: begin
				q			<=			16'hD91F;
		end
		32'h00005764: begin
				q			<=			16'h2083;
		end
		32'h00005766: begin
				q			<=			16'h00C1;
		end
		32'h00005768: begin
				q			<=			16'h3513;
		end
		32'h0000576A: begin
				q			<=			16'h0015;
		end
		32'h0000576C: begin
				q			<=			16'h0113;
		end
		32'h0000576E: begin
				q			<=			16'h0101;
		end
		32'h00005770: begin
				q			<=			16'h8067;
		end
		32'h00005772: begin
				q			<=			16'h0000;
		end
		32'h00005774: begin
				q			<=			16'h0513;
		end
		32'h00005776: begin
				q			<=			16'h0000;
		end
		32'h00005778: begin
				q			<=			16'h8067;
		end
		32'h0000577A: begin
				q			<=			16'h0000;
		end
		32'h0000577C: begin
				q			<=			16'h0793;
		end
		32'h0000577E: begin
				q			<=			16'h0125;
		end
		32'h00005780: begin
				q			<=			16'h0513;
		end
		32'h00005782: begin
				q			<=			16'h0025;
		end
		32'h00005784: begin
				q			<=			16'h1F23;
		end
		32'h00005786: begin
				q			<=			16'hFE05;
		end
		32'h00005788: begin
				q			<=			16'h1CE3;
		end
		32'h0000578A: begin
				q			<=			16'hFEF5;
		end
		32'h0000578C: begin
				q			<=			16'h5783;
		end
		32'h0000578E: begin
				q			<=			16'h0005;
		end
		32'h00005790: begin
				q			<=			16'h8737;
		end
		32'h00005792: begin
				q			<=			16'h0000;
		end
		32'h00005794: begin
				q			<=			16'h0713;
		end
		32'h00005796: begin
				q			<=			16'hFFF7;
		end
		32'h00005798: begin
				q			<=			16'hE7B3;
		end
		32'h0000579A: begin
				q			<=			16'h00E7;
		end
		32'h0000579C: begin
				q			<=			16'h1023;
		end
		32'h0000579E: begin
				q			<=			16'h00F5;
		end
		32'h000057A0: begin
				q			<=			16'h8067;
		end
		32'h000057A2: begin
				q			<=			16'h0000;
		end
		32'h000057A4: begin
				q			<=			16'h0113;
		end
		32'h000057A6: begin
				q			<=			16'hFE01;
		end
		32'h000057A8: begin
				q			<=			16'h2C23;
		end
		32'h000057AA: begin
				q			<=			16'h0081;
		end
		32'h000057AC: begin
				q			<=			16'h2623;
		end
		32'h000057AE: begin
				q			<=			16'h0131;
		end
		32'h000057B0: begin
				q			<=			16'h2E23;
		end
		32'h000057B2: begin
				q			<=			16'h0011;
		end
		32'h000057B4: begin
				q			<=			16'h2A23;
		end
		32'h000057B6: begin
				q			<=			16'h0091;
		end
		32'h000057B8: begin
				q			<=			16'h2823;
		end
		32'h000057BA: begin
				q			<=			16'h0121;
		end
		32'h000057BC: begin
				q			<=			16'h2423;
		end
		32'h000057BE: begin
				q			<=			16'h0141;
		end
		32'h000057C0: begin
				q			<=			16'h2223;
		end
		32'h000057C2: begin
				q			<=			16'h0151;
		end
		32'h000057C4: begin
				q			<=			16'h0993;
		end
		32'h000057C6: begin
				q			<=			16'h0005;
		end
		32'h000057C8: begin
				q			<=			16'h8413;
		end
		32'h000057CA: begin
				q			<=			16'h0005;
		end
		32'h000057CC: begin
				q			<=			16'hD863;
		end
		32'h000057CE: begin
				q			<=			16'h1005;
		end
		32'h000057D0: begin
				q			<=			16'h0933;
		end
		32'h000057D2: begin
				q			<=			16'h40B0;
		end
		32'h000057D4: begin
				q			<=			16'h0A13;
		end
		32'h000057D6: begin
				q			<=			16'h0009;
		end
		32'h000057D8: begin
				q			<=			16'h0493;
		end
		32'h000057DA: begin
				q			<=			16'h0000;
		end
		32'h000057DC: begin
				q			<=			16'h0A93;
		end
		32'h000057DE: begin
				q			<=			16'h00F0;
		end
		32'h000057E0: begin
				q			<=			16'hCE63;
		end
		32'h000057E2: begin
				q			<=			16'h034A;
		end
		32'h000057E4: begin
				q			<=			16'h5913;
		end
		32'h000057E6: begin
				q			<=			16'h0049;
		end
		32'h000057E8: begin
				q			<=			16'h0593;
		end
		32'h000057EA: begin
				q			<=			16'hFF00;
		end
		32'h000057EC: begin
				q			<=			16'h05B3;
		end
		32'h000057EE: begin
				q			<=			16'h02B9;
		end
		32'h000057F0: begin
				q			<=			16'h0A13;
		end
		32'h000057F2: begin
				q			<=			16'h0070;
		end
		32'h000057F4: begin
				q			<=			16'h8433;
		end
		32'h000057F6: begin
				q			<=			16'h4085;
		end
		32'h000057F8: begin
				q			<=			16'h0913;
		end
		32'h000057FA: begin
				q			<=			16'h0004;
		end
		32'h000057FC: begin
				q			<=			16'h4C63;
		end
		32'h000057FE: begin
				q			<=			16'h032A;
		end
		32'h00005800: begin
				q			<=			16'h5593;
		end
		32'h00005802: begin
				q			<=			16'h0034;
		end
		32'h00005804: begin
				q			<=			16'h0793;
		end
		32'h00005806: begin
				q			<=			16'hFF80;
		end
		32'h00005808: begin
				q			<=			16'h85B3;
		end
		32'h0000580A: begin
				q			<=			16'h02F5;
		end
		32'h0000580C: begin
				q			<=			16'h8433;
		end
		32'h0000580E: begin
				q			<=			16'h0085;
		end
		32'h00005810: begin
				q			<=			16'h1063;
		end
		32'h00005812: begin
				q			<=			16'h0404;
		end
		32'h00005814: begin
				q			<=			16'h3533;
		end
		32'h00005816: begin
				q			<=			16'h0090;
		end
		32'h00005818: begin
				q			<=			16'h006F;
		end
		32'h0000581A: begin
				q			<=			16'h0A00;
		end
		32'h0000581C: begin
				q			<=			16'hD783;
		end
		32'h0000581E: begin
				q			<=			16'h0189;
		end
		32'h00005820: begin
				q			<=			16'h8513;
		end
		32'h00005822: begin
				q			<=			16'h0009;
		end
		32'h00005824: begin
				q			<=			16'h0A13;
		end
		32'h00005826: begin
				q			<=			16'hFF0A;
		end
		32'h00005828: begin
				q			<=			16'hE4B3;
		end
		32'h0000582A: begin
				q			<=			16'h00F4;
		end
		32'h0000582C: begin
				q			<=			16'hF0EF;
		end
		32'h0000582E: begin
				q			<=			16'hB91F;
		end
		32'h00005830: begin
				q			<=			16'hF06F;
		end
		32'h00005832: begin
				q			<=			16'hFB1F;
		end
		32'h00005834: begin
				q			<=			16'hC783;
		end
		32'h00005836: begin
				q			<=			16'h0189;
		end
		32'h00005838: begin
				q			<=			16'h8513;
		end
		32'h0000583A: begin
				q			<=			16'h0009;
		end
		32'h0000583C: begin
				q			<=			16'h0913;
		end
		32'h0000583E: begin
				q			<=			16'hFF89;
		end
		32'h00005840: begin
				q			<=			16'hE4B3;
		end
		32'h00005842: begin
				q			<=			16'h0097;
		end
		32'h00005844: begin
				q			<=			16'h0097;
		end
		32'h00005846: begin
				q			<=			16'h0000;
		end
		32'h00005848: begin
				q			<=			16'h80E7;
		end
		32'h0000584A: begin
				q			<=			16'hAFC0;
		end
		32'h0000584C: begin
				q			<=			16'hF06F;
		end
		32'h0000584E: begin
				q			<=			16'hFB1F;
		end
		32'h00005850: begin
				q			<=			16'hD783;
		end
		32'h00005852: begin
				q			<=			16'h0189;
		end
		32'h00005854: begin
				q			<=			16'h8513;
		end
		32'h00005856: begin
				q			<=			16'h0009;
		end
		32'h00005858: begin
				q			<=			16'h0413;
		end
		32'h0000585A: begin
				q			<=			16'hFFF4;
		end
		32'h0000585C: begin
				q			<=			16'hF793;
		end
		32'h0000585E: begin
				q			<=			16'h0017;
		end
		32'h00005860: begin
				q			<=			16'hE4B3;
		end
		32'h00005862: begin
				q			<=			16'h0097;
		end
		32'h00005864: begin
				q			<=			16'h0097;
		end
		32'h00005866: begin
				q			<=			16'h0000;
		end
		32'h00005868: begin
				q			<=			16'h80E7;
		end
		32'h0000586A: begin
				q			<=			16'hA380;
		end
		32'h0000586C: begin
				q			<=			16'hF06F;
		end
		32'h0000586E: begin
				q			<=			16'hFA5F;
		end
		32'h00005870: begin
				q			<=			16'h8513;
		end
		32'h00005872: begin
				q			<=			16'h0009;
		end
		32'h00005874: begin
				q			<=			16'h0097;
		end
		32'h00005876: begin
				q			<=			16'h0000;
		end
		32'h00005878: begin
				q			<=			16'h80E7;
		end
		32'h0000587A: begin
				q			<=			16'hB280;
		end
		32'h0000587C: begin
				q			<=			16'h8493;
		end
		32'h0000587E: begin
				q			<=			16'hFF04;
		end
		32'h00005880: begin
				q			<=			16'h48E3;
		end
		32'h00005882: begin
				q			<=			16'hFE99;
		end
		32'h00005884: begin
				q			<=			16'h5593;
		end
		32'h00005886: begin
				q			<=			16'h0044;
		end
		32'h00005888: begin
				q			<=			16'h0793;
		end
		32'h0000588A: begin
				q			<=			16'hFF00;
		end
		32'h0000588C: begin
				q			<=			16'h85B3;
		end
		32'h0000588E: begin
				q			<=			16'h02F5;
		end
		32'h00005890: begin
				q			<=			16'h0913;
		end
		32'h00005892: begin
				q			<=			16'h0070;
		end
		32'h00005894: begin
				q			<=			16'h0433;
		end
		32'h00005896: begin
				q			<=			16'h00B4;
		end
		32'h00005898: begin
				q			<=			16'h0493;
		end
		32'h0000589A: begin
				q			<=			16'h0004;
		end
		32'h0000589C: begin
				q			<=			16'h4663;
		end
		32'h0000589E: begin
				q			<=			16'h0499;
		end
		32'h000058A0: begin
				q			<=			16'h5593;
		end
		32'h000058A2: begin
				q			<=			16'h0034;
		end
		32'h000058A4: begin
				q			<=			16'h0793;
		end
		32'h000058A6: begin
				q			<=			16'hFF80;
		end
		32'h000058A8: begin
				q			<=			16'h85B3;
		end
		32'h000058AA: begin
				q			<=			16'h02F5;
		end
		32'h000058AC: begin
				q			<=			16'h0433;
		end
		32'h000058AE: begin
				q			<=			16'h00B4;
		end
		32'h000058B0: begin
				q			<=			16'h1463;
		end
		32'h000058B2: begin
				q			<=			16'h0404;
		end
		32'h000058B4: begin
				q			<=			16'h0513;
		end
		32'h000058B6: begin
				q			<=			16'h0000;
		end
		32'h000058B8: begin
				q			<=			16'h2083;
		end
		32'h000058BA: begin
				q			<=			16'h01C1;
		end
		32'h000058BC: begin
				q			<=			16'h2403;
		end
		32'h000058BE: begin
				q			<=			16'h0181;
		end
		32'h000058C0: begin
				q			<=			16'h2483;
		end
		32'h000058C2: begin
				q			<=			16'h0141;
		end
		32'h000058C4: begin
				q			<=			16'h2903;
		end
		32'h000058C6: begin
				q			<=			16'h0101;
		end
		32'h000058C8: begin
				q			<=			16'h2983;
		end
		32'h000058CA: begin
				q			<=			16'h00C1;
		end
		32'h000058CC: begin
				q			<=			16'h2A03;
		end
		32'h000058CE: begin
				q			<=			16'h0081;
		end
		32'h000058D0: begin
				q			<=			16'h2A83;
		end
		32'h000058D2: begin
				q			<=			16'h0041;
		end
		32'h000058D4: begin
				q			<=			16'h0113;
		end
		32'h000058D6: begin
				q			<=			16'h0201;
		end
		32'h000058D8: begin
				q			<=			16'h8067;
		end
		32'h000058DA: begin
				q			<=			16'h0000;
		end
		32'h000058DC: begin
				q			<=			16'h8493;
		end
		32'h000058DE: begin
				q			<=			16'h0005;
		end
		32'h000058E0: begin
				q			<=			16'h0913;
		end
		32'h000058E2: begin
				q			<=			16'h00F0;
		end
		32'h000058E4: begin
				q			<=			16'hF06F;
		end
		32'h000058E6: begin
				q			<=			16'hF9DF;
		end
		32'h000058E8: begin
				q			<=			16'h8513;
		end
		32'h000058EA: begin
				q			<=			16'h0009;
		end
		32'h000058EC: begin
				q			<=			16'hF0EF;
		end
		32'h000058EE: begin
				q			<=			16'hA89F;
		end
		32'h000058F0: begin
				q			<=			16'h8493;
		end
		32'h000058F2: begin
				q			<=			16'hFF84;
		end
		32'h000058F4: begin
				q			<=			16'hF06F;
		end
		32'h000058F6: begin
				q			<=			16'hFA9F;
		end
		32'h000058F8: begin
				q			<=			16'h8513;
		end
		32'h000058FA: begin
				q			<=			16'h0009;
		end
		32'h000058FC: begin
				q			<=			16'hF0EF;
		end
		32'h000058FE: begin
				q			<=			16'h9F1F;
		end
		32'h00005900: begin
				q			<=			16'h0413;
		end
		32'h00005902: begin
				q			<=			16'hFFF4;
		end
		32'h00005904: begin
				q			<=			16'hF06F;
		end
		32'h00005906: begin
				q			<=			16'hFADF;
		end
		32'h00005908: begin
				q			<=			16'h5783;
		end
		32'h0000590A: begin
				q			<=			16'h0045;
		end
		32'h0000590C: begin
				q			<=			16'h0113;
		end
		32'h0000590E: begin
				q			<=			16'hFF01;
		end
		32'h00005910: begin
				q			<=			16'h2223;
		end
		32'h00005912: begin
				q			<=			16'h0091;
		end
		32'h00005914: begin
				q			<=			16'h2623;
		end
		32'h00005916: begin
				q			<=			16'h0011;
		end
		32'h00005918: begin
				q			<=			16'h2423;
		end
		32'h0000591A: begin
				q			<=			16'h0081;
		end
		32'h0000591C: begin
				q			<=			16'h2023;
		end
		32'h0000591E: begin
				q			<=			16'h0121;
		end
		32'h00005920: begin
				q			<=			16'h0493;
		end
		32'h00005922: begin
				q			<=			16'h0005;
		end
		32'h00005924: begin
				q			<=			16'h9663;
		end
		32'h00005926: begin
				q			<=			16'h0807;
		end
		32'h00005928: begin
				q			<=			16'h1783;
		end
		32'h0000592A: begin
				q			<=			16'h0065;
		end
		32'h0000592C: begin
				q			<=			16'h0413;
		end
		32'h0000592E: begin
				q			<=			16'h0000;
		end
		32'h00005930: begin
				q			<=			16'h0913;
		end
		32'h00005932: begin
				q			<=			16'h0A00;
		end
		32'h00005934: begin
				q			<=			16'hD863;
		end
		32'h00005936: begin
				q			<=			16'h0207;
		end
		32'h00005938: begin
				q			<=			16'h0513;
		end
		32'h0000593A: begin
				q			<=			16'h0004;
		end
		32'h0000593C: begin
				q			<=			16'h2083;
		end
		32'h0000593E: begin
				q			<=			16'h00C1;
		end
		32'h00005940: begin
				q			<=			16'h2403;
		end
		32'h00005942: begin
				q			<=			16'h0081;
		end
		32'h00005944: begin
				q			<=			16'h2483;
		end
		32'h00005946: begin
				q			<=			16'h0041;
		end
		32'h00005948: begin
				q			<=			16'h2903;
		end
		32'h0000594A: begin
				q			<=			16'h0001;
		end
		32'h0000594C: begin
				q			<=			16'h0113;
		end
		32'h0000594E: begin
				q			<=			16'h0101;
		end
		32'h00005950: begin
				q			<=			16'h8067;
		end
		32'h00005952: begin
				q			<=			16'h0000;
		end
		32'h00005954: begin
				q			<=			16'h8513;
		end
		32'h00005956: begin
				q			<=			16'h0004;
		end
		32'h00005958: begin
				q			<=			16'h0413;
		end
		32'h0000595A: begin
				q			<=			16'h0104;
		end
		32'h0000595C: begin
				q			<=			16'hF0EF;
		end
		32'h0000595E: begin
				q			<=			16'hA41F;
		end
		32'h00005960: begin
				q			<=			16'h0CE3;
		end
		32'h00005962: begin
				q			<=			16'hFD24;
		end
		32'h00005964: begin
				q			<=			16'hD783;
		end
		32'h00005966: begin
				q			<=			16'h0064;
		end
		32'h00005968: begin
				q			<=			16'h86E3;
		end
		32'h0000596A: begin
				q			<=			16'hFE07;
		end
		32'h0000596C: begin
				q			<=			16'hD783;
		end
		32'h0000596E: begin
				q			<=			16'h0064;
		end
		32'h00005970: begin
				q			<=			16'hF793;
		end
		32'h00005972: begin
				q			<=			16'hF007;
		end
		32'h00005974: begin
				q			<=			16'h8463;
		end
		32'h00005976: begin
				q			<=			16'h0207;
		end
		32'h00005978: begin
				q			<=			16'h0913;
		end
		32'h0000597A: begin
				q			<=			16'h0A00;
		end
		32'h0000597C: begin
				q			<=			16'h9783;
		end
		32'h0000597E: begin
				q			<=			16'h0064;
		end
		32'h00005980: begin
				q			<=			16'hCCE3;
		end
		32'h00005982: begin
				q			<=			16'hFA07;
		end
		32'h00005984: begin
				q			<=			16'h8513;
		end
		32'h00005986: begin
				q			<=			16'h0004;
		end
		32'h00005988: begin
				q			<=			16'h0413;
		end
		32'h0000598A: begin
				q			<=			16'h0014;
		end
		32'h0000598C: begin
				q			<=			16'h0097;
		end
		32'h0000598E: begin
				q			<=			16'h0000;
		end
		32'h00005990: begin
				q			<=			16'h80E7;
		end
		32'h00005992: begin
				q			<=			16'h9600;
		end
		32'h00005994: begin
				q			<=			16'h54E3;
		end
		32'h00005996: begin
				q			<=			16'hFE89;
		end
		32'h00005998: begin
				q			<=			16'hF06F;
		end
		32'h0000599A: begin
				q			<=			16'hFA1F;
		end
		32'h0000599C: begin
				q			<=			16'h8513;
		end
		32'h0000599E: begin
				q			<=			16'h0004;
		end
		32'h000059A0: begin
				q			<=			16'h0097;
		end
		32'h000059A2: begin
				q			<=			16'h0000;
		end
		32'h000059A4: begin
				q			<=			16'h80E7;
		end
		32'h000059A6: begin
				q			<=			16'h9D40;
		end
		32'h000059A8: begin
				q			<=			16'h0413;
		end
		32'h000059AA: begin
				q			<=			16'h0084;
		end
		32'h000059AC: begin
				q			<=			16'hF06F;
		end
		32'h000059AE: begin
				q			<=			16'hFC1F;
		end
		32'h000059B0: begin
				q			<=			16'hF793;
		end
		32'h000059B2: begin
				q			<=			16'hF007;
		end
		32'h000059B4: begin
				q			<=			16'h0413;
		end
		32'h000059B6: begin
				q			<=			16'h0000;
		end
		32'h000059B8: begin
				q			<=			16'h8663;
		end
		32'h000059BA: begin
				q			<=			16'h0007;
		end
		32'h000059BC: begin
				q			<=			16'hF0EF;
		end
		32'h000059BE: begin
				q			<=			16'h985F;
		end
		32'h000059C0: begin
				q			<=			16'h0413;
		end
		32'h000059C2: begin
				q			<=			16'hFF80;
		end
		32'h000059C4: begin
				q			<=			16'h0913;
		end
		32'h000059C6: begin
				q			<=			16'hF700;
		end
		32'h000059C8: begin
				q			<=			16'h006F;
		end
		32'h000059CA: begin
				q			<=			16'h0140;
		end
		32'h000059CC: begin
				q			<=			16'h8513;
		end
		32'h000059CE: begin
				q			<=			16'h0004;
		end
		32'h000059D0: begin
				q			<=			16'h0413;
		end
		32'h000059D2: begin
				q			<=			16'hFFF4;
		end
		32'h000059D4: begin
				q			<=			16'hF0EF;
		end
		32'h000059D6: begin
				q			<=			16'h8C9F;
		end
		32'h000059D8: begin
				q			<=			16'h40E3;
		end
		32'h000059DA: begin
				q			<=			16'hF724;
		end
		32'h000059DC: begin
				q			<=			16'hD783;
		end
		32'h000059DE: begin
				q			<=			16'h0044;
		end
		32'h000059E0: begin
				q			<=			16'h96E3;
		end
		32'h000059E2: begin
				q			<=			16'hFE07;
		end
		32'h000059E4: begin
				q			<=			16'hF06F;
		end
		32'h000059E6: begin
				q			<=			16'hF55F;
		end
		32'h000059E8: begin
				q			<=			16'h0793;
		end
		32'h000059EA: begin
				q			<=			16'h0105;
		end
		32'h000059EC: begin
				q			<=			16'h0513;
		end
		32'h000059EE: begin
				q			<=			16'h0025;
		end
		32'h000059F0: begin
				q			<=			16'h1F23;
		end
		32'h000059F2: begin
				q			<=			16'hFE05;
		end
		32'h000059F4: begin
				q			<=			16'h1CE3;
		end
		32'h000059F6: begin
				q			<=			16'hFEF5;
		end
		32'h000059F8: begin
				q			<=			16'hC7B7;
		end
		32'h000059FA: begin
				q			<=			16'hFFFF;
		end
		32'h000059FC: begin
				q			<=			16'h1023;
		end
		32'h000059FE: begin
				q			<=			16'h00F5;
		end
		32'h00005A00: begin
				q			<=			16'h87B7;
		end
		32'h00005A02: begin
				q			<=			16'h0000;
		end
		32'h00005A04: begin
				q			<=			16'h8793;
		end
		32'h00005A06: begin
				q			<=			16'hFFF7;
		end
		32'h00005A08: begin
				q			<=			16'h1123;
		end
		32'h00005A0A: begin
				q			<=			16'h00F5;
		end
		32'h00005A0C: begin
				q			<=			16'h8067;
		end
		32'h00005A0E: begin
				q			<=			16'h0000;
		end
		32'h00005A10: begin
				q			<=			16'h0713;
		end
		32'h00005A12: begin
				q			<=			16'h0005;
		end
		32'h00005A14: begin
				q			<=			16'h5683;
		end
		32'h00005A16: begin
				q			<=			16'h0007;
		end
		32'h00005A18: begin
				q			<=			16'h8513;
		end
		32'h00005A1A: begin
				q			<=			16'h0005;
		end
		32'h00005A1C: begin
				q			<=			16'h5783;
		end
		32'h00005A1E: begin
				q			<=			16'h0027;
		end
		32'h00005A20: begin
				q			<=			16'h8663;
		end
		32'h00005A22: begin
				q			<=			16'h0006;
		end
		32'h00005A24: begin
				q			<=			16'h86B7;
		end
		32'h00005A26: begin
				q			<=			16'hFFFF;
		end
		32'h00005A28: begin
				q			<=			16'hE7B3;
		end
		32'h00005A2A: begin
				q			<=			16'h00D7;
		end
		32'h00005A2C: begin
				q			<=			16'h1923;
		end
		32'h00005A2E: begin
				q			<=			16'h00F5;
		end
		32'h00005A30: begin
				q			<=			16'h5603;
		end
		32'h00005A32: begin
				q			<=			16'h0027;
		end
		32'h00005A34: begin
				q			<=			16'h86B7;
		end
		32'h00005A36: begin
				q			<=			16'h0000;
		end
		32'h00005A38: begin
				q			<=			16'h8693;
		end
		32'h00005A3A: begin
				q			<=			16'hFFF6;
		end
		32'h00005A3C: begin
				q			<=			16'h0793;
		end
		32'h00005A3E: begin
				q			<=			16'h0067;
		end
		32'h00005A40: begin
				q			<=			16'h1E63;
		end
		32'h00005A42: begin
				q			<=			16'h00D6;
		end
		32'h00005A44: begin
				q			<=			16'h0713;
		end
		32'h00005A46: begin
				q			<=			16'h01A7;
		end
		32'h00005A48: begin
				q			<=			16'hD683;
		end
		32'h00005A4A: begin
				q			<=			16'h0007;
		end
		32'h00005A4C: begin
				q			<=			16'h9863;
		end
		32'h00005A4E: begin
				q			<=			16'h0206;
		end
		32'h00005A50: begin
				q			<=			16'h8793;
		end
		32'h00005A52: begin
				q			<=			16'h0027;
		end
		32'h00005A54: begin
				q			<=			16'h9AE3;
		end
		32'h00005A56: begin
				q			<=			16'hFEE7;
		end
		32'h00005A58: begin
				q			<=			16'hF06F;
		end
		32'h00005A5A: begin
				q			<=			16'hD25F;
		end
		32'h00005A5C: begin
				q			<=			16'h0513;
		end
		32'h00005A5E: begin
				q			<=			16'h0105;
		end
		32'h00005A60: begin
				q			<=			16'h0713;
		end
		32'h00005A62: begin
				q			<=			16'h0187;
		end
		32'h00005A64: begin
				q			<=			16'h8793;
		end
		32'h00005A66: begin
				q			<=			16'h0027;
		end
		32'h00005A68: begin
				q			<=			16'hD683;
		end
		32'h00005A6A: begin
				q			<=			16'hFFE7;
		end
		32'h00005A6C: begin
				q			<=			16'h0513;
		end
		32'h00005A6E: begin
				q			<=			16'hFFE5;
		end
		32'h00005A70: begin
				q			<=			16'h1123;
		end
		32'h00005A72: begin
				q			<=			16'h00D5;
		end
		32'h00005A74: begin
				q			<=			16'h98E3;
		end
		32'h00005A76: begin
				q			<=			16'hFEE7;
		end
		32'h00005A78: begin
				q			<=			16'h8067;
		end
		32'h00005A7A: begin
				q			<=			16'h0000;
		end
		32'h00005A7C: begin
				q			<=			16'h0317;
		end
		32'h00005A7E: begin
				q			<=			16'h0000;
		end
		32'h00005A80: begin
				q			<=			16'h0067;
		end
		32'h00005A82: begin
				q			<=			16'hF6C3;
		end
		32'h00005A84: begin
				q			<=			16'h0113;
		end
		32'h00005A86: begin
				q			<=			16'hFD01;
		end
		32'h00005A88: begin
				q			<=			16'h2223;
		end
		32'h00005A8A: begin
				q			<=			16'h0291;
		end
		32'h00005A8C: begin
				q			<=			16'h0493;
		end
		32'h00005A8E: begin
				q			<=			16'h0005;
		end
		32'h00005A90: begin
				q			<=			16'h0513;
		end
		32'h00005A92: begin
				q			<=			16'h0041;
		end
		32'h00005A94: begin
				q			<=			16'h2423;
		end
		32'h00005A96: begin
				q			<=			16'h0281;
		end
		32'h00005A98: begin
				q			<=			16'h2623;
		end
		32'h00005A9A: begin
				q			<=			16'h0211;
		end
		32'h00005A9C: begin
				q			<=			16'h8413;
		end
		32'h00005A9E: begin
				q			<=			16'h0005;
		end
		32'h00005AA0: begin
				q			<=			16'hF0EF;
		end
		32'h00005AA2: begin
				q			<=			16'hF88F;
		end
		32'h00005AA4: begin
				q			<=			16'hD703;
		end
		32'h00005AA6: begin
				q			<=			16'h00E4;
		end
		32'h00005AA8: begin
				q			<=			16'h1793;
		end
		32'h00005AAA: begin
				q			<=			16'h0107;
		end
		32'h00005AAC: begin
				q			<=			16'hD793;
		end
		32'h00005AAE: begin
				q			<=			16'h4107;
		end
		32'h00005AB0: begin
				q			<=			16'hC263;
		end
		32'h00005AB2: begin
				q			<=			16'h0407;
		end
		32'h00005AB4: begin
				q			<=			16'h1223;
		end
		32'h00005AB6: begin
				q			<=			16'h0001;
		end
		32'h00005AB8: begin
				q			<=			16'h86B7;
		end
		32'h00005ABA: begin
				q			<=			16'h0000;
		end
		32'h00005ABC: begin
				q			<=			16'h8693;
		end
		32'h00005ABE: begin
				q			<=			16'hFFF6;
		end
		32'h00005AC0: begin
				q			<=			16'h7733;
		end
		32'h00005AC2: begin
				q			<=			16'h00D7;
		end
		32'h00005AC4: begin
				q			<=			16'h8793;
		end
		32'h00005AC6: begin
				q			<=			16'h00E4;
		end
		32'h00005AC8: begin
				q			<=			16'h1E63;
		end
		32'h00005ACA: begin
				q			<=			16'h06D7;
		end
		32'h00005ACC: begin
				q			<=			16'h8713;
		end
		32'h00005ACE: begin
				q			<=			16'h0004;
		end
		32'h00005AD0: begin
				q			<=			16'h5683;
		end
		32'h00005AD2: begin
				q			<=			16'h0007;
		end
		32'h00005AD4: begin
				q			<=			16'h8663;
		end
		32'h00005AD6: begin
				q			<=			16'h0206;
		end
		32'h00005AD8: begin
				q			<=			16'h0513;
		end
		32'h00005ADA: begin
				q			<=			16'h0004;
		end
		32'h00005ADC: begin
				q			<=			16'hF0EF;
		end
		32'h00005ADE: begin
				q			<=			16'hF0DF;
		end
		32'h00005AE0: begin
				q			<=			16'h2083;
		end
		32'h00005AE2: begin
				q			<=			16'h02C1;
		end
		32'h00005AE4: begin
				q			<=			16'h2403;
		end
		32'h00005AE6: begin
				q			<=			16'h0281;
		end
		32'h00005AE8: begin
				q			<=			16'h2483;
		end
		32'h00005AEA: begin
				q			<=			16'h0241;
		end
		32'h00005AEC: begin
				q			<=			16'h0113;
		end
		32'h00005AEE: begin
				q			<=			16'h0301;
		end
		32'h00005AF0: begin
				q			<=			16'h8067;
		end
		32'h00005AF2: begin
				q			<=			16'h0000;
		end
		32'h00005AF4: begin
				q			<=			16'h0793;
		end
		32'h00005AF6: begin
				q			<=			16'hFFF0;
		end
		32'h00005AF8: begin
				q			<=			16'h1223;
		end
		32'h00005AFA: begin
				q			<=			16'h00F1;
		end
		32'h00005AFC: begin
				q			<=			16'hF06F;
		end
		32'h00005AFE: begin
				q			<=			16'hFBDF;
		end
		32'h00005B00: begin
				q			<=			16'h0713;
		end
		32'h00005B02: begin
				q			<=			16'h0027;
		end
		32'h00005B04: begin
				q			<=			16'h96E3;
		end
		32'h00005B06: begin
				q			<=			16'hFCE7;
		end
		32'h00005B08: begin
				q			<=			16'h0513;
		end
		32'h00005B0A: begin
				q			<=			16'h0004;
		end
		32'h00005B0C: begin
				q			<=			16'hF0EF;
		end
		32'h00005B0E: begin
				q			<=			16'hEECF;
		end
		32'h00005B10: begin
				q			<=			16'h0513;
		end
		32'h00005B12: begin
				q			<=			16'h0004;
		end
		32'h00005B14: begin
				q			<=			16'h0097;
		end
		32'h00005B16: begin
				q			<=			16'h0000;
		end
		32'h00005B18: begin
				q			<=			16'h80E7;
		end
		32'h00005B1A: begin
				q			<=			16'hC680;
		end
		32'h00005B1C: begin
				q			<=			16'h9783;
		end
		32'h00005B1E: begin
				q			<=			16'h00E4;
		end
		32'h00005B20: begin
				q			<=			16'hD0E3;
		end
		32'h00005B22: begin
				q			<=			16'hFC07;
		end
		32'h00005B24: begin
				q			<=			16'h0513;
		end
		32'h00005B26: begin
				q			<=			16'h0004;
		end
		32'h00005B28: begin
				q			<=			16'hF0EF;
		end
		32'h00005B2A: begin
				q			<=			16'h9C9F;
		end
		32'h00005B2C: begin
				q			<=			16'h1AE3;
		end
		32'h00005B2E: begin
				q			<=			16'hFA05;
		end
		32'h00005B30: begin
				q			<=			16'h5783;
		end
		32'h00005B32: begin
				q			<=			16'h0124;
		end
		32'h00005B34: begin
				q			<=			16'h8737;
		end
		32'h00005B36: begin
				q			<=			16'hFFFF;
		end
		32'h00005B38: begin
				q			<=			16'hC7B3;
		end
		32'h00005B3A: begin
				q			<=			16'h00E7;
		end
		32'h00005B3C: begin
				q			<=			16'h1923;
		end
		32'h00005B3E: begin
				q			<=			16'h00F4;
		end
		32'h00005B40: begin
				q			<=			16'hF06F;
		end
		32'h00005B42: begin
				q			<=			16'hFA1F;
		end
		32'h00005B44: begin
				q			<=			16'h1323;
		end
		32'h00005B46: begin
				q			<=			16'h00E1;
		end
		32'h00005B48: begin
				q			<=			16'h0693;
		end
		32'h00005B4A: begin
				q			<=			16'h0041;
		end
		32'h00005B4C: begin
				q			<=			16'h8793;
		end
		32'h00005B4E: begin
				q			<=			16'hFFE7;
		end
		32'h00005B50: begin
				q			<=			16'hD603;
		end
		32'h00005B52: begin
				q			<=			16'h0007;
		end
		32'h00005B54: begin
				q			<=			16'h8693;
		end
		32'h00005B56: begin
				q			<=			16'h0026;
		end
		32'h00005B58: begin
				q			<=			16'h9223;
		end
		32'h00005B5A: begin
				q			<=			16'h00C6;
		end
		32'h00005B5C: begin
				q			<=			16'h98E3;
		end
		32'h00005B5E: begin
				q			<=			16'hFEF4;
		end
		32'h00005B60: begin
				q			<=			16'h1E63;
		end
		32'h00005B62: begin
				q			<=			16'h0007;
		end
		32'h00005B64: begin
				q			<=			16'h1423;
		end
		32'h00005B66: begin
				q			<=			16'h0001;
		end
		32'h00005B68: begin
				q			<=			16'h0593;
		end
		32'h00005B6A: begin
				q			<=			16'h0004;
		end
		32'h00005B6C: begin
				q			<=			16'h0513;
		end
		32'h00005B6E: begin
				q			<=			16'h0041;
		end
		32'h00005B70: begin
				q			<=			16'h0097;
		end
		32'h00005B72: begin
				q			<=			16'h0000;
		end
		32'h00005B74: begin
				q			<=			16'h80E7;
		end
		32'h00005B76: begin
				q			<=			16'hEA00;
		end
		32'h00005B78: begin
				q			<=			16'hF06F;
		end
		32'h00005B7A: begin
				q			<=			16'hF69F;
		end
		32'h00005B7C: begin
				q			<=			16'h0793;
		end
		32'h00005B7E: begin
				q			<=			16'h0010;
		end
		32'h00005B80: begin
				q			<=			16'h0593;
		end
		32'h00005B82: begin
				q			<=			16'hFFF0;
		end
		32'h00005B84: begin
				q			<=			16'h0513;
		end
		32'h00005B86: begin
				q			<=			16'h0041;
		end
		32'h00005B88: begin
				q			<=			16'h1423;
		end
		32'h00005B8A: begin
				q			<=			16'h00F1;
		end
		32'h00005B8C: begin
				q			<=			16'hF0EF;
		end
		32'h00005B8E: begin
				q			<=			16'hC19F;
		end
		32'h00005B90: begin
				q			<=			16'hF06F;
		end
		32'h00005B92: begin
				q			<=			16'hFD9F;
		end
		32'h00005B94: begin
				q			<=			16'h0113;
		end
		32'h00005B96: begin
				q			<=			16'hFE01;
		end
		32'h00005B98: begin
				q			<=			16'h2C23;
		end
		32'h00005B9A: begin
				q			<=			16'h0081;
		end
		32'h00005B9C: begin
				q			<=			16'h2A23;
		end
		32'h00005B9E: begin
				q			<=			16'h0091;
		end
		32'h00005BA0: begin
				q			<=			16'h2823;
		end
		32'h00005BA2: begin
				q			<=			16'h0121;
		end
		32'h00005BA4: begin
				q			<=			16'h2623;
		end
		32'h00005BA6: begin
				q			<=			16'h0131;
		end
		32'h00005BA8: begin
				q			<=			16'h2423;
		end
		32'h00005BAA: begin
				q			<=			16'h0141;
		end
		32'h00005BAC: begin
				q			<=			16'h2223;
		end
		32'h00005BAE: begin
				q			<=			16'h0151;
		end
		32'h00005BB0: begin
				q			<=			16'h8913;
		end
		32'h00005BB2: begin
				q			<=			16'h0006;
		end
		32'h00005BB4: begin
				q			<=			16'h8413;
		end
		32'h00005BB6: begin
				q			<=			16'h0007;
		end
		32'h00005BB8: begin
				q			<=			16'h2E23;
		end
		32'h00005BBA: begin
				q			<=			16'h0011;
		end
		32'h00005BBC: begin
				q			<=			16'h0493;
		end
		32'h00005BBE: begin
				q			<=			16'h0005;
		end
		32'h00005BC0: begin
				q			<=			16'h8993;
		end
		32'h00005BC2: begin
				q			<=			16'h0005;
		end
		32'h00005BC4: begin
				q			<=			16'h0A13;
		end
		32'h00005BC6: begin
				q			<=			16'h0006;
		end
		32'h00005BC8: begin
				q			<=			16'h0A93;
		end
		32'h00005BCA: begin
				q			<=			16'h0007;
		end
		32'h00005BCC: begin
				q			<=			16'hF0EF;
		end
		32'h00005BCE: begin
				q			<=			16'hD3DF;
		end
		32'h00005BD0: begin
				q			<=			16'h0793;
		end
		32'h00005BD2: begin
				q			<=			16'h0900;
		end
		32'h00005BD4: begin
				q			<=			16'h0933;
		end
		32'h00005BD6: begin
				q			<=			16'h40A9;
		end
		32'h00005BD8: begin
				q			<=			16'hD463;
		end
		32'h00005BDA: begin
				q			<=			16'h04A7;
		end
		32'h00005BDC: begin
				q			<=			16'h87B7;
		end
		32'h00005BDE: begin
				q			<=			16'h0000;
		end
		32'h00005BE0: begin
				q			<=			16'h8793;
		end
		32'h00005BE2: begin
				q			<=			16'hFFE7;
		end
		32'h00005BE4: begin
				q			<=			16'hCC63;
		end
		32'h00005BE6: begin
				q			<=			16'h2D27;
		end
		32'h00005BE8: begin
				q			<=			16'h8793;
		end
		32'h00005BEA: begin
				q			<=			16'h0024;
		end
		32'h00005BEC: begin
				q			<=			16'h8493;
		end
		32'h00005BEE: begin
				q			<=			16'h01A4;
		end
		32'h00005BF0: begin
				q			<=			16'h8793;
		end
		32'h00005BF2: begin
				q			<=			16'h0027;
		end
		32'h00005BF4: begin
				q			<=			16'h9F23;
		end
		32'h00005BF6: begin
				q			<=			16'hFE07;
		end
		32'h00005BF8: begin
				q			<=			16'h9CE3;
		end
		32'h00005BFA: begin
				q			<=			16'hFE97;
		end
		32'h00005BFC: begin
				q			<=			16'h2083;
		end
		32'h00005BFE: begin
				q			<=			16'h01C1;
		end
		32'h00005C00: begin
				q			<=			16'h2403;
		end
		32'h00005C02: begin
				q			<=			16'h0181;
		end
		32'h00005C04: begin
				q			<=			16'h2483;
		end
		32'h00005C06: begin
				q			<=			16'h0141;
		end
		32'h00005C08: begin
				q			<=			16'h2903;
		end
		32'h00005C0A: begin
				q			<=			16'h0101;
		end
		32'h00005C0C: begin
				q			<=			16'h2983;
		end
		32'h00005C0E: begin
				q			<=			16'h00C1;
		end
		32'h00005C10: begin
				q			<=			16'h2A03;
		end
		32'h00005C12: begin
				q			<=			16'h0081;
		end
		32'h00005C14: begin
				q			<=			16'h2A83;
		end
		32'h00005C16: begin
				q			<=			16'h0041;
		end
		32'h00005C18: begin
				q			<=			16'h0113;
		end
		32'h00005C1A: begin
				q			<=			16'h0201;
		end
		32'h00005C1C: begin
				q			<=			16'h8067;
		end
		32'h00005C1E: begin
				q			<=			16'h0000;
		end
		32'h00005C20: begin
				q			<=			16'h5063;
		end
		32'h00005C22: begin
				q			<=			16'h0209;
		end
		32'h00005C24: begin
				q			<=			16'h0793;
		end
		32'h00005C26: begin
				q			<=			16'hF700;
		end
		32'h00005C28: begin
				q			<=			16'h4063;
		end
		32'h00005C2A: begin
				q			<=			16'h14F9;
		end
		32'h00005C2C: begin
				q			<=			16'h0593;
		end
		32'h00005C2E: begin
				q			<=			16'h0009;
		end
		32'h00005C30: begin
				q			<=			16'h8513;
		end
		32'h00005C32: begin
				q			<=			16'h0004;
		end
		32'h00005C34: begin
				q			<=			16'h0097;
		end
		32'h00005C36: begin
				q			<=			16'h0000;
		end
		32'h00005C38: begin
				q			<=			16'h80E7;
		end
		32'h00005C3A: begin
				q			<=			16'hB700;
		end
		32'h00005C3C: begin
				q			<=			16'h1263;
		end
		32'h00005C3E: begin
				q			<=			16'h1405;
		end
		32'h00005C40: begin
				q			<=			16'h8A63;
		end
		32'h00005C42: begin
				q			<=			16'h220A;
		end
		32'h00005C44: begin
				q			<=			16'h2703;
		end
		32'h00005C46: begin
				q			<=			16'h0044;
		end
		32'h00005C48: begin
				q			<=			16'h2783;
		end
		32'h00005C4A: begin
				q			<=			16'h0004;
		end
		32'h00005C4C: begin
				q			<=			16'h0863;
		end
		32'h00005C4E: begin
				q			<=			16'h06F7;
		end
		32'h00005C50: begin
				q			<=			16'h0513;
		end
		32'h00005C52: begin
				q			<=			16'h01A4;
		end
		32'h00005C54: begin
				q			<=			16'hF097;
		end
		32'h00005C56: begin
				q			<=			16'hFFFF;
		end
		32'h00005C58: begin
				q			<=			16'h80E7;
		end
		32'h00005C5A: begin
				q			<=			16'h5D40;
		end
		32'h00005C5C: begin
				q			<=			16'h2783;
		end
		32'h00005C5E: begin
				q			<=			16'h0044;
		end
		32'h00005C60: begin
				q			<=			16'h0713;
		end
		32'h00005C62: begin
				q			<=			16'h0380;
		end
		32'h00005C64: begin
				q			<=			16'h8E63;
		end
		32'h00005C66: begin
				q			<=			16'h16E7;
		end
		32'h00005C68: begin
				q			<=			16'h4063;
		end
		32'h00005C6A: begin
				q			<=			16'h12F7;
		end
		32'h00005C6C: begin
				q			<=			16'h0713;
		end
		32'h00005C6E: begin
				q			<=			16'h0180;
		end
		32'h00005C70: begin
				q			<=			16'h8663;
		end
		32'h00005C72: begin
				q			<=			16'h1AE7;
		end
		32'h00005C74: begin
				q			<=			16'h0713;
		end
		32'h00005C76: begin
				q			<=			16'h0350;
		end
		32'h00005C78: begin
				q			<=			16'h8263;
		end
		32'h00005C7A: begin
				q			<=			16'h18E7;
		end
		32'h00005C7C: begin
				q			<=			16'h0713;
		end
		32'h00005C7E: begin
				q			<=			16'h00C0;
		end
		32'h00005C80: begin
				q			<=			16'h2423;
		end
		32'h00005C82: begin
				q			<=			16'h00E4;
		end
		32'h00005C84: begin
				q			<=			16'h0737;
		end
		32'h00005C86: begin
				q			<=			16'h8001;
		end
		32'h00005C88: begin
				q			<=			16'h0713;
		end
		32'h00005C8A: begin
				q			<=			16'hFFF7;
		end
		32'h00005C8C: begin
				q			<=			16'h2A23;
		end
		32'h00005C8E: begin
				q			<=			16'h00E4;
		end
		32'h00005C90: begin
				q			<=			16'h0713;
		end
		32'h00005C92: begin
				q			<=			16'h0010;
		end
		32'h00005C94: begin
				q			<=			16'h1C23;
		end
		32'h00005C96: begin
				q			<=			16'h00E4;
		end
		32'h00005C98: begin
				q			<=			16'h0713;
		end
		32'h00005C9A: begin
				q			<=			16'h00B0;
		end
		32'h00005C9C: begin
				q			<=			16'h2623;
		end
		32'h00005C9E: begin
				q			<=			16'h00E4;
		end
		32'h00005CA0: begin
				q			<=			16'h2703;
		end
		32'h00005CA2: begin
				q			<=			16'h00C4;
		end
		32'h00005CA4: begin
				q			<=			16'h5683;
		end
		32'h00005CA6: begin
				q			<=			16'h0184;
		end
		32'h00005CA8: begin
				q			<=			16'h0713;
		end
		32'h00005CAA: begin
				q			<=			16'h0087;
		end
		32'h00005CAC: begin
				q			<=			16'h1713;
		end
		32'h00005CAE: begin
				q			<=			16'h0017;
		end
		32'h00005CB0: begin
				q			<=			16'h0733;
		end
		32'h00005CB2: begin
				q			<=			16'h00E4;
		end
		32'h00005CB4: begin
				q			<=			16'h1523;
		end
		32'h00005CB6: begin
				q			<=			16'h00D7;
		end
		32'h00005CB8: begin
				q			<=			16'h2023;
		end
		32'h00005CBA: begin
				q			<=			16'h00F4;
		end
		32'h00005CBC: begin
				q			<=			16'h4263;
		end
		32'h00005CBE: begin
				q			<=			16'h0320;
		end
		32'h00005CC0: begin
				q			<=			16'h2703;
		end
		32'h00005CC2: begin
				q			<=			16'h0044;
		end
		32'h00005CC4: begin
				q			<=			16'h0793;
		end
		32'h00005CC6: begin
				q			<=			16'h0900;
		end
		32'h00005CC8: begin
				q			<=			16'h0C63;
		end
		32'h00005CCA: begin
				q			<=			16'h00F7;
		end
		32'h00005CCC: begin
				q			<=			16'hD783;
		end
		32'h00005CCE: begin
				q			<=			16'h0184;
		end
		32'h00005CD0: begin
				q			<=			16'h8513;
		end
		32'h00005CD2: begin
				q			<=			16'h0004;
		end
		32'h00005CD4: begin
				q			<=			16'hF793;
		end
		32'h00005CD6: begin
				q			<=			16'h0017;
		end
		32'h00005CD8: begin
				q			<=			16'hE9B3;
		end
		32'h00005CDA: begin
				q			<=			16'h00F9;
		end
		32'h00005CDC: begin
				q			<=			16'hF0EF;
		end
		32'h00005CDE: begin
				q			<=			16'hDC0F;
		end
		32'h00005CE0: begin
				q			<=			16'h2683;
		end
		32'h00005CE2: begin
				q			<=			16'h0084;
		end
		32'h00005CE4: begin
				q			<=			16'h5603;
		end
		32'h00005CE6: begin
				q			<=			16'h0144;
		end
		32'h00005CE8: begin
				q			<=			16'h2583;
		end
		32'h00005CEA: begin
				q			<=			16'h0044;
		end
		32'h00005CEC: begin
				q			<=			16'h9713;
		end
		32'h00005CEE: begin
				q			<=			16'h0016;
		end
		32'h00005CF0: begin
				q			<=			16'h8733;
		end
		32'h00005CF2: begin
				q			<=			16'h00E4;
		end
		32'h00005CF4: begin
				q			<=			16'h5783;
		end
		32'h00005CF6: begin
				q			<=			16'h0007;
		end
		32'h00005CF8: begin
				q			<=			16'hF7B3;
		end
		32'h00005CFA: begin
				q			<=			16'h00C7;
		end
		32'h00005CFC: begin
				q			<=			16'h0613;
		end
		32'h00005CFE: begin
				q			<=			16'h08F0;
		end
		32'h00005D00: begin
				q			<=			16'h4A63;
		end
		32'h00005D02: begin
				q			<=			16'h00B6;
		end
		32'h00005D04: begin
				q			<=			16'h8693;
		end
		32'h00005D06: begin
				q			<=			16'h0016;
		end
		32'h00005D08: begin
				q			<=			16'h0613;
		end
		32'h00005D0A: begin
				q			<=			16'h0007;
		end
		32'h00005D0C: begin
				q			<=			16'h0593;
		end
		32'h00005D0E: begin
				q			<=			16'h00C0;
		end
		32'h00005D10: begin
				q			<=			16'hDA63;
		end
		32'h00005D12: begin
				q			<=			16'h10D5;
		end
		32'h00005D14: begin
				q			<=			16'h5683;
		end
		32'h00005D16: begin
				q			<=			16'h0144;
		end
		32'h00005D18: begin
				q			<=			16'h5603;
		end
		32'h00005D1A: begin
				q			<=			16'h0007;
		end
		32'h00005D1C: begin
				q			<=			16'hC693;
		end
		32'h00005D1E: begin
				q			<=			16'hFFF6;
		end
		32'h00005D20: begin
				q			<=			16'hF6B3;
		end
		32'h00005D22: begin
				q			<=			16'h00C6;
		end
		32'h00005D24: begin
				q			<=			16'h1023;
		end
		32'h00005D26: begin
				q			<=			16'h00D7;
		end
		32'h00005D28: begin
				q			<=			16'h5703;
		end
		32'h00005D2A: begin
				q			<=			16'h0164;
		end
		32'h00005D2C: begin
				q			<=			16'h76B3;
		end
		32'h00005D2E: begin
				q			<=			16'h00F7;
		end
		32'h00005D30: begin
				q			<=			16'h8A63;
		end
		32'h00005D32: begin
				q			<=			16'h1006;
		end
		32'h00005D34: begin
				q			<=			16'h1263;
		end
		32'h00005D36: begin
				q			<=			16'h02F7;
		end
		32'h00005D38: begin
				q			<=			16'h9463;
		end
		32'h00005D3A: begin
				q			<=			16'h1009;
		end
		32'h00005D3C: begin
				q			<=			16'h2783;
		end
		32'h00005D3E: begin
				q			<=			16'h00C4;
		end
		32'h00005D40: begin
				q			<=			16'h5703;
		end
		32'h00005D42: begin
				q			<=			16'h0184;
		end
		32'h00005D44: begin
				q			<=			16'h9793;
		end
		32'h00005D46: begin
				q			<=			16'h0017;
		end
		32'h00005D48: begin
				q			<=			16'h87B3;
		end
		32'h00005D4A: begin
				q			<=			16'h00F4;
		end
		32'h00005D4C: begin
				q			<=			16'hD783;
		end
		32'h00005D4E: begin
				q			<=			16'h0007;
		end
		32'h00005D50: begin
				q			<=			16'hF7B3;
		end
		32'h00005D52: begin
				q			<=			16'h00E7;
		end
		32'h00005D54: begin
				q			<=			16'h8863;
		end
		32'h00005D56: begin
				q			<=			16'h0E07;
		end
		32'h00005D58: begin
				q			<=			16'h8593;
		end
		32'h00005D5A: begin
				q			<=			16'h0004;
		end
		32'h00005D5C: begin
				q			<=			16'h0513;
		end
		32'h00005D5E: begin
				q			<=			16'h01A4;
		end
		32'h00005D60: begin
				q			<=			16'hF0EF;
		end
		32'h00005D62: begin
				q			<=			16'hE84F;
		end
		32'h00005D64: begin
				q			<=			16'h006F;
		end
		32'h00005D66: begin
				q			<=			16'h0E00;
		end
		32'h00005D68: begin
				q			<=			16'h8793;
		end
		32'h00005D6A: begin
				q			<=			16'h0024;
		end
		32'h00005D6C: begin
				q			<=			16'h8493;
		end
		32'h00005D6E: begin
				q			<=			16'h01A4;
		end
		32'h00005D70: begin
				q			<=			16'h8793;
		end
		32'h00005D72: begin
				q			<=			16'h0027;
		end
		32'h00005D74: begin
				q			<=			16'h9F23;
		end
		32'h00005D76: begin
				q			<=			16'hFE07;
		end
		32'h00005D78: begin
				q			<=			16'h9CE3;
		end
		32'h00005D7A: begin
				q			<=			16'hFE97;
		end
		32'h00005D7C: begin
				q			<=			16'hF06F;
		end
		32'h00005D7E: begin
				q			<=			16'hE81F;
		end
		32'h00005D80: begin
				q			<=			16'h0993;
		end
		32'h00005D82: begin
				q			<=			16'h0010;
		end
		32'h00005D84: begin
				q			<=			16'hF06F;
		end
		32'h00005D86: begin
				q			<=			16'hEBDF;
		end
		32'h00005D88: begin
				q			<=			16'h0713;
		end
		32'h00005D8A: begin
				q			<=			16'h0400;
		end
		32'h00005D8C: begin
				q			<=			16'h8863;
		end
		32'h00005D8E: begin
				q			<=			16'h02E7;
		end
		32'h00005D90: begin
				q			<=			16'h0713;
		end
		32'h00005D92: begin
				q			<=			16'h0710;
		end
		32'h00005D94: begin
				q			<=			16'h94E3;
		end
		32'h00005D96: begin
				q			<=			16'hEEE7;
		end
		32'h00005D98: begin
				q			<=			16'h8737;
		end
		32'h00005D9A: begin
				q			<=			16'h4000;
		end
		32'h00005D9C: begin
				q			<=			16'h0713;
		end
		32'h00005D9E: begin
				q			<=			16'hFFF7;
		end
		32'h00005DA0: begin
				q			<=			16'h0693;
		end
		32'h00005DA2: begin
				q			<=			16'h00A0;
		end
		32'h00005DA4: begin
				q			<=			16'h2A23;
		end
		32'h00005DA6: begin
				q			<=			16'h00E4;
		end
		32'h00005DA8: begin
				q			<=			16'h2423;
		end
		32'h00005DAA: begin
				q			<=			16'h00D4;
		end
		32'h00005DAC: begin
				q			<=			16'h8737;
		end
		32'h00005DAE: begin
				q			<=			16'hFFFF;
		end
		32'h00005DB0: begin
				q			<=			16'h1C23;
		end
		32'h00005DB2: begin
				q			<=			16'h00E4;
		end
		32'h00005DB4: begin
				q			<=			16'h2623;
		end
		32'h00005DB6: begin
				q			<=			16'h00D4;
		end
		32'h00005DB8: begin
				q			<=			16'hF06F;
		end
		32'h00005DBA: begin
				q			<=			16'hEE9F;
		end
		32'h00005DBC: begin
				q			<=			16'h0713;
		end
		32'h00005DBE: begin
				q			<=			16'h0070;
		end
		32'h00005DC0: begin
				q			<=			16'h2423;
		end
		32'h00005DC2: begin
				q			<=			16'h00E4;
		end
		32'h00005DC4: begin
				q			<=			16'h0737;
		end
		32'h00005DC6: begin
				q			<=			16'h8001;
		end
		32'h00005DC8: begin
				q			<=			16'h0713;
		end
		32'h00005DCA: begin
				q			<=			16'hFFF7;
		end
		32'h00005DCC: begin
				q			<=			16'h2A23;
		end
		32'h00005DCE: begin
				q			<=			16'h00E4;
		end
		32'h00005DD0: begin
				q			<=			16'h0713;
		end
		32'h00005DD2: begin
				q			<=			16'h0010;
		end
		32'h00005DD4: begin
				q			<=			16'h1C23;
		end
		32'h00005DD6: begin
				q			<=			16'h00E4;
		end
		32'h00005DD8: begin
				q			<=			16'h0713;
		end
		32'h00005DDA: begin
				q			<=			16'h0060;
		end
		32'h00005DDC: begin
				q			<=			16'hF06F;
		end
		32'h00005DDE: begin
				q			<=			16'hEC1F;
		end
		32'h00005DE0: begin
				q			<=			16'h0693;
		end
		32'h00005DE2: begin
				q			<=			16'h0060;
		end
		32'h00005DE4: begin
				q			<=			16'h0737;
		end
		32'h00005DE6: begin
				q			<=			16'h0080;
		end
		32'h00005DE8: begin
				q			<=			16'h0713;
		end
		32'h00005DEA: begin
				q			<=			16'h0FF7;
		end
		32'h00005DEC: begin
				q			<=			16'h2A23;
		end
		32'h00005DEE: begin
				q			<=			16'h00E4;
		end
		32'h00005DF0: begin
				q			<=			16'h2423;
		end
		32'h00005DF2: begin
				q			<=			16'h00D4;
		end
		32'h00005DF4: begin
				q			<=			16'h0713;
		end
		32'h00005DF6: begin
				q			<=			16'h1000;
		end
		32'h00005DF8: begin
				q			<=			16'hF06F;
		end
		32'h00005DFA: begin
				q			<=			16'hFB9F;
		end
		32'h00005DFC: begin
				q			<=			16'h0737;
		end
		32'h00005DFE: begin
				q			<=			16'h0400;
		end
		32'h00005E00: begin
				q			<=			16'h0713;
		end
		32'h00005E02: begin
				q			<=			16'h7FF7;
		end
		32'h00005E04: begin
				q			<=			16'h0693;
		end
		32'h00005E06: begin
				q			<=			16'h0060;
		end
		32'h00005E08: begin
				q			<=			16'h2A23;
		end
		32'h00005E0A: begin
				q			<=			16'h00E4;
		end
		32'h00005E0C: begin
				q			<=			16'h1737;
		end
		32'h00005E0E: begin
				q			<=			16'h0000;
		end
		32'h00005E10: begin
				q			<=			16'h2423;
		end
		32'h00005E12: begin
				q			<=			16'h00D4;
		end
		32'h00005E14: begin
				q			<=			16'h0713;
		end
		32'h00005E16: begin
				q			<=			16'h8007;
		end
		32'h00005E18: begin
				q			<=			16'hF06F;
		end
		32'h00005E1A: begin
				q			<=			16'hF99F;
		end
		32'h00005E1C: begin
				q			<=			16'h0693;
		end
		32'h00005E1E: begin
				q			<=			16'h0040;
		end
		32'h00005E20: begin
				q			<=			16'hF06F;
		end
		32'h00005E22: begin
				q			<=			16'hFC5F;
		end
		32'h00005E24: begin
				q			<=			16'h5503;
		end
		32'h00005E26: begin
				q			<=			16'h0026;
		end
		32'h00005E28: begin
				q			<=			16'h0463;
		end
		32'h00005E2A: begin
				q			<=			16'h0005;
		end
		32'h00005E2C: begin
				q			<=			16'hE793;
		end
		32'h00005E2E: begin
				q			<=			16'h0017;
		end
		32'h00005E30: begin
				q			<=			16'h1123;
		end
		32'h00005E32: begin
				q			<=			16'h0006;
		end
		32'h00005E34: begin
				q			<=			16'h8693;
		end
		32'h00005E36: begin
				q			<=			16'h0016;
		end
		32'h00005E38: begin
				q			<=			16'h0613;
		end
		32'h00005E3A: begin
				q			<=			16'h0026;
		end
		32'h00005E3C: begin
				q			<=			16'hF06F;
		end
		32'h00005E3E: begin
				q			<=			16'hED5F;
		end
		32'h00005E40: begin
				q			<=			16'h0CE3;
		end
		32'h00005E42: begin
				q			<=			16'hF00A;
		end
		32'h00005E44: begin
				q			<=			16'h4E63;
		end
		32'h00005E46: begin
				q			<=			16'h0120;
		end
		32'h00005E48: begin
				q			<=			16'h2703;
		end
		32'h00005E4A: begin
				q			<=			16'h0044;
		end
		32'h00005E4C: begin
				q			<=			16'h0793;
		end
		32'h00005E4E: begin
				q			<=			16'h0900;
		end
		32'h00005E50: begin
				q			<=			16'h0863;
		end
		32'h00005E52: begin
				q			<=			16'h00F7;
		end
		32'h00005E54: begin
				q			<=			16'h8513;
		end
		32'h00005E56: begin
				q			<=			16'h0004;
		end
		32'h00005E58: begin
				q			<=			16'hF097;
		end
		32'h00005E5A: begin
				q			<=			16'hFFFF;
		end
		32'h00005E5C: begin
				q			<=			16'h80E7;
		end
		32'h00005E5E: begin
				q			<=			16'h4940;
		end
		32'h00005E60: begin
				q			<=			16'hD783;
		end
		32'h00005E62: begin
				q			<=			16'h0044;
		end
		32'h00005E64: begin
				q			<=			16'h8863;
		end
		32'h00005E66: begin
				q			<=			16'h0007;
		end
		32'h00005E68: begin
				q			<=			16'h8513;
		end
		32'h00005E6A: begin
				q			<=			16'h0004;
		end
		32'h00005E6C: begin
				q			<=			16'hF0EF;
		end
		32'h00005E6E: begin
				q			<=			16'hC30F;
		end
		32'h00005E70: begin
				q			<=			16'h0913;
		end
		32'h00005E72: begin
				q			<=			16'h0019;
		end
		32'h00005E74: begin
				q			<=			16'h87B7;
		end
		32'h00005E76: begin
				q			<=			16'h0000;
		end
		32'h00005E78: begin
				q			<=			16'h9C23;
		end
		32'h00005E7A: begin
				q			<=			16'h0004;
		end
		32'h00005E7C: begin
				q			<=			16'h8793;
		end
		32'h00005E7E: begin
				q			<=			16'hFFE7;
		end
		32'h00005E80: begin
				q			<=			16'hD463;
		end
		32'h00005E82: begin
				q			<=			16'h0327;
		end
		32'h00005E84: begin
				q			<=			16'h87B7;
		end
		32'h00005E86: begin
				q			<=			16'hFFFF;
		end
		32'h00005E88: begin
				q			<=			16'hC793;
		end
		32'h00005E8A: begin
				q			<=			16'hFFF7;
		end
		32'h00005E8C: begin
				q			<=			16'h9123;
		end
		32'h00005E8E: begin
				q			<=			16'h00F4;
		end
		32'h00005E90: begin
				q			<=			16'h8793;
		end
		32'h00005E92: begin
				q			<=			16'h0044;
		end
		32'h00005E94: begin
				q			<=			16'h8493;
		end
		32'h00005E96: begin
				q			<=			16'h0184;
		end
		32'h00005E98: begin
				q			<=			16'h9023;
		end
		32'h00005E9A: begin
				q			<=			16'h0007;
		end
		32'h00005E9C: begin
				q			<=			16'h8793;
		end
		32'h00005E9E: begin
				q			<=			16'h0027;
		end
		32'h00005EA0: begin
				q			<=			16'h9CE3;
		end
		32'h00005EA2: begin
				q			<=			16'hFEF4;
		end
		32'h00005EA4: begin
				q			<=			16'hF06F;
		end
		32'h00005EA6: begin
				q			<=			16'hD59F;
		end
		32'h00005EA8: begin
				q			<=			16'h5663;
		end
		32'h00005EAA: begin
				q			<=			16'h0009;
		end
		32'h00005EAC: begin
				q			<=			16'h9123;
		end
		32'h00005EAE: begin
				q			<=			16'h0004;
		end
		32'h00005EB0: begin
				q			<=			16'hF06F;
		end
		32'h00005EB2: begin
				q			<=			16'hD4DF;
		end
		32'h00005EB4: begin
				q			<=			16'h9123;
		end
		32'h00005EB6: begin
				q			<=			16'h0124;
		end
		32'h00005EB8: begin
				q			<=			16'hF06F;
		end
		32'h00005EBA: begin
				q			<=			16'hD45F;
		end
		32'h00005EBC: begin
				q			<=			16'h94E3;
		end
		32'h00005EBE: begin
				q			<=			16'hD80A;
		end
		32'h00005EC0: begin
				q			<=			16'h9C23;
		end
		32'h00005EC2: begin
				q			<=			16'h0004;
		end
		32'h00005EC4: begin
				q			<=			16'hF06F;
		end
		32'h00005EC6: begin
				q			<=			16'hFC1F;
		end
		32'h00005EC8: begin
				q			<=			16'h0113;
		end
		32'h00005ECA: begin
				q			<=			16'hFE01;
		end
		32'h00005ECC: begin
				q			<=			16'h2423;
		end
		32'h00005ECE: begin
				q			<=			16'h0141;
		end
		32'h00005ED0: begin
				q			<=			16'h5A03;
		end
		32'h00005ED2: begin
				q			<=			16'h0025;
		end
		32'h00005ED4: begin
				q			<=			16'h2C23;
		end
		32'h00005ED6: begin
				q			<=			16'h0081;
		end
		32'h00005ED8: begin
				q			<=			16'h8413;
		end
		32'h00005EDA: begin
				q			<=			16'h0005;
		end
		32'h00005EDC: begin
				q			<=			16'h2E23;
		end
		32'h00005EDE: begin
				q			<=			16'h0011;
		end
		32'h00005EE0: begin
				q			<=			16'h2A23;
		end
		32'h00005EE2: begin
				q			<=			16'h0091;
		end
		32'h00005EE4: begin
				q			<=			16'h2823;
		end
		32'h00005EE6: begin
				q			<=			16'h0121;
		end
		32'h00005EE8: begin
				q			<=			16'h2223;
		end
		32'h00005EEA: begin
				q			<=			16'h0151;
		end
		32'h00005EEC: begin
				q			<=			16'h2023;
		end
		32'h00005EEE: begin
				q			<=			16'h0161;
		end
		32'h00005EF0: begin
				q			<=			16'h0913;
		end
		32'h00005EF2: begin
				q			<=			16'h0006;
		end
		32'h00005EF4: begin
				q			<=			16'h0B13;
		end
		32'h00005EF6: begin
				q			<=			16'h0346;
		end
		32'h00005EF8: begin
				q			<=			16'h2623;
		end
		32'h00005EFA: begin
				q			<=			16'h0131;
		end
		32'h00005EFC: begin
				q			<=			16'h0A93;
		end
		32'h00005EFE: begin
				q			<=			16'h0005;
		end
		32'h00005F00: begin
				q			<=			16'h0097;
		end
		32'h00005F02: begin
				q			<=			16'h0000;
		end
		32'h00005F04: begin
				q			<=			16'h80E7;
		end
		32'h00005F06: begin
				q			<=			16'hA080;
		end
		32'h00005F08: begin
				q			<=			16'h5483;
		end
		32'h00005F0A: begin
				q			<=			16'h0024;
		end
		32'h00005F0C: begin
				q			<=			16'h0A33;
		end
		32'h00005F0E: begin
				q			<=			16'h40AA;
		end
		32'h00005F10: begin
				q			<=			16'h0513;
		end
		32'h00005F12: begin
				q			<=			16'h0004;
		end
		32'h00005F14: begin
				q			<=			16'h0097;
		end
		32'h00005F16: begin
				q			<=			16'h0000;
		end
		32'h00005F18: begin
				q			<=			16'h80E7;
		end
		32'h00005F1A: begin
				q			<=			16'h9F40;
		end
		32'h00005F1C: begin
				q			<=			16'h84B3;
		end
		32'h00005F1E: begin
				q			<=			16'h40A4;
		end
		32'h00005F20: begin
				q			<=			16'h0513;
		end
		32'h00005F22: begin
				q			<=			16'h000B;
		end
		32'h00005F24: begin
				q			<=			16'hF0EF;
		end
		32'h00005F26: begin
				q			<=			16'hB04F;
		end
		32'h00005F28: begin
				q			<=			16'hD463;
		end
		32'h00005F2A: begin
				q			<=			16'h0544;
		end
		32'h00005F2C: begin
				q			<=			16'h0513;
		end
		32'h00005F2E: begin
				q			<=			16'h0004;
		end
		32'h00005F30: begin
				q			<=			16'h2403;
		end
		32'h00005F32: begin
				q			<=			16'h0181;
		end
		32'h00005F34: begin
				q			<=			16'h2083;
		end
		32'h00005F36: begin
				q			<=			16'h01C1;
		end
		32'h00005F38: begin
				q			<=			16'h2983;
		end
		32'h00005F3A: begin
				q			<=			16'h00C1;
		end
		32'h00005F3C: begin
				q			<=			16'h2A03;
		end
		32'h00005F3E: begin
				q			<=			16'h0081;
		end
		32'h00005F40: begin
				q			<=			16'h2A83;
		end
		32'h00005F42: begin
				q			<=			16'h0041;
		end
		32'h00005F44: begin
				q			<=			16'h2B03;
		end
		32'h00005F46: begin
				q			<=			16'h0001;
		end
		32'h00005F48: begin
				q			<=			16'h0793;
		end
		32'h00005F4A: begin
				q			<=			16'h0009;
		end
		32'h00005F4C: begin
				q			<=			16'h8693;
		end
		32'h00005F4E: begin
				q			<=			16'h0004;
		end
		32'h00005F50: begin
				q			<=			16'h2903;
		end
		32'h00005F52: begin
				q			<=			16'h0101;
		end
		32'h00005F54: begin
				q			<=			16'h2483;
		end
		32'h00005F56: begin
				q			<=			16'h0141;
		end
		32'h00005F58: begin
				q			<=			16'h0713;
		end
		32'h00005F5A: begin
				q			<=			16'h0000;
		end
		32'h00005F5C: begin
				q			<=			16'h0613;
		end
		32'h00005F5E: begin
				q			<=			16'h0000;
		end
		32'h00005F60: begin
				q			<=			16'h0593;
		end
		32'h00005F62: begin
				q			<=			16'h0000;
		end
		32'h00005F64: begin
				q			<=			16'h0113;
		end
		32'h00005F66: begin
				q			<=			16'h0201;
		end
		32'h00005F68: begin
				q			<=			16'h0317;
		end
		32'h00005F6A: begin
				q			<=			16'h0000;
		end
		32'h00005F6C: begin
				q			<=			16'h0067;
		end
		32'h00005F6E: begin
				q			<=			16'hC2C3;
		end
		32'h00005F70: begin
				q			<=			16'h0593;
		end
		32'h00005F72: begin
				q			<=			16'h0004;
		end
		32'h00005F74: begin
				q			<=			16'h8513;
		end
		32'h00005F76: begin
				q			<=			16'h000A;
		end
		32'h00005F78: begin
				q			<=			16'hF0EF;
		end
		32'h00005F7A: begin
				q			<=			16'hAE8F;
		end
		32'h00005F7C: begin
				q			<=			16'h0993;
		end
		32'h00005F7E: begin
				q			<=			16'h0000;
		end
		32'h00005F80: begin
				q			<=			16'h4A63;
		end
		32'h00005F82: begin
				q			<=			16'h00A0;
		end
		32'h00005F84: begin
				q			<=			16'h0593;
		end
		32'h00005F86: begin
				q			<=			16'h0004;
		end
		32'h00005F88: begin
				q			<=			16'h8513;
		end
		32'h00005F8A: begin
				q			<=			16'h000A;
		end
		32'h00005F8C: begin
				q			<=			16'hF0EF;
		end
		32'h00005F8E: begin
				q			<=			16'hC90F;
		end
		32'h00005F90: begin
				q			<=			16'h0993;
		end
		32'h00005F92: begin
				q			<=			16'h0010;
		end
		32'h00005F94: begin
				q			<=			16'h0513;
		end
		32'h00005F96: begin
				q			<=			16'h000B;
		end
		32'h00005F98: begin
				q			<=			16'hF0EF;
		end
		32'h00005F9A: begin
				q			<=			16'hB54F;
		end
		32'h00005F9C: begin
				q			<=			16'h5783;
		end
		32'h00005F9E: begin
				q			<=			16'h04C9;
		end
		32'h00005FA0: begin
				q			<=			16'h0513;
		end
		32'h00005FA2: begin
				q			<=			16'h0004;
		end
		32'h00005FA4: begin
				q			<=			16'h8493;
		end
		32'h00005FA6: begin
				q			<=			16'hFFF4;
		end
		32'h00005FA8: begin
				q			<=			16'hE9B3;
		end
		32'h00005FAA: begin
				q			<=			16'h00F9;
		end
		32'h00005FAC: begin
				q			<=			16'h1623;
		end
		32'h00005FAE: begin
				q			<=			16'h0539;
		end
		32'h00005FB0: begin
				q			<=			16'hF0EF;
		end
		32'h00005FB2: begin
				q			<=			16'hB3CF;
		end
		32'h00005FB4: begin
				q			<=			16'hF06F;
		end
		32'h00005FB6: begin
				q			<=			16'hF75F;
		end
		32'h00005FB8: begin
				q			<=			16'h0113;
		end
		32'h00005FBA: begin
				q			<=			16'hF701;
		end
		32'h00005FBC: begin
				q			<=			16'h2423;
		end
		32'h00005FBE: begin
				q			<=			16'h0881;
		end
		32'h00005FC0: begin
				q			<=			16'h2223;
		end
		32'h00005FC2: begin
				q			<=			16'h0891;
		end
		32'h00005FC4: begin
				q			<=			16'h2023;
		end
		32'h00005FC6: begin
				q			<=			16'h0921;
		end
		32'h00005FC8: begin
				q			<=			16'h2E23;
		end
		32'h00005FCA: begin
				q			<=			16'h0731;
		end
		32'h00005FCC: begin
				q			<=			16'h2623;
		end
		32'h00005FCE: begin
				q			<=			16'h0811;
		end
		32'h00005FD0: begin
				q			<=			16'h2C23;
		end
		32'h00005FD2: begin
				q			<=			16'h0741;
		end
		32'h00005FD4: begin
				q			<=			16'h2A23;
		end
		32'h00005FD6: begin
				q			<=			16'h0751;
		end
		32'h00005FD8: begin
				q			<=			16'h2823;
		end
		32'h00005FDA: begin
				q			<=			16'h0761;
		end
		32'h00005FDC: begin
				q			<=			16'h2623;
		end
		32'h00005FDE: begin
				q			<=			16'h0771;
		end
		32'h00005FE0: begin
				q			<=			16'h2423;
		end
		32'h00005FE2: begin
				q			<=			16'h0781;
		end
		32'h00005FE4: begin
				q			<=			16'h2223;
		end
		32'h00005FE6: begin
				q			<=			16'h0791;
		end
		32'h00005FE8: begin
				q			<=			16'h0493;
		end
		32'h00005FEA: begin
				q			<=			16'h0005;
		end
		32'h00005FEC: begin
				q			<=			16'h8413;
		end
		32'h00005FEE: begin
				q			<=			16'h0005;
		end
		32'h00005FF0: begin
				q			<=			16'h0913;
		end
		32'h00005FF2: begin
				q			<=			16'h0006;
		end
		32'h00005FF4: begin
				q			<=			16'h8993;
		end
		32'h00005FF6: begin
				q			<=			16'h0006;
		end
		32'h00005FF8: begin
				q			<=			16'hF097;
		end
		32'h00005FFA: begin
				q			<=			16'hFFFF;
		end
		32'h00005FFC: begin
				q			<=			16'h80E7;
		end
		32'h00005FFE: begin
				q			<=			16'h4F80;
		end
		32'h00006000: begin
				q			<=			16'h0263;
		end
		32'h00006002: begin
				q			<=			16'h0405;
		end
		32'h00006004: begin
				q			<=			16'h0593;
		end
		32'h00006006: begin
				q			<=			16'h0009;
		end
		32'h00006008: begin
				q			<=			16'h8513;
		end
		32'h0000600A: begin
				q			<=			16'h0004;
		end
		32'h0000600C: begin
				q			<=			16'hF0EF;
		end
		32'h0000600E: begin
				q			<=			16'hA00F;
		end
		32'h00006010: begin
				q			<=			16'h2083;
		end
		32'h00006012: begin
				q			<=			16'h08C1;
		end
		32'h00006014: begin
				q			<=			16'h2403;
		end
		32'h00006016: begin
				q			<=			16'h0881;
		end
		32'h00006018: begin
				q			<=			16'h2483;
		end
		32'h0000601A: begin
				q			<=			16'h0841;
		end
		32'h0000601C: begin
				q			<=			16'h2903;
		end
		32'h0000601E: begin
				q			<=			16'h0801;
		end
		32'h00006020: begin
				q			<=			16'h2983;
		end
		32'h00006022: begin
				q			<=			16'h07C1;
		end
		32'h00006024: begin
				q			<=			16'h2A03;
		end
		32'h00006026: begin
				q			<=			16'h0781;
		end
		32'h00006028: begin
				q			<=			16'h2A83;
		end
		32'h0000602A: begin
				q			<=			16'h0741;
		end
		32'h0000602C: begin
				q			<=			16'h2B03;
		end
		32'h0000602E: begin
				q			<=			16'h0701;
		end
		32'h00006030: begin
				q			<=			16'h2B83;
		end
		32'h00006032: begin
				q			<=			16'h06C1;
		end
		32'h00006034: begin
				q			<=			16'h2C03;
		end
		32'h00006036: begin
				q			<=			16'h0681;
		end
		32'h00006038: begin
				q			<=			16'h2C83;
		end
		32'h0000603A: begin
				q			<=			16'h0641;
		end
		32'h0000603C: begin
				q			<=			16'h0113;
		end
		32'h0000603E: begin
				q			<=			16'h0901;
		end
		32'h00006040: begin
				q			<=			16'h8067;
		end
		32'h00006042: begin
				q			<=			16'h0000;
		end
		32'h00006044: begin
				q			<=			16'h0513;
		end
		32'h00006046: begin
				q			<=			16'h0004;
		end
		32'h00006048: begin
				q			<=			16'hF097;
		end
		32'h0000604A: begin
				q			<=			16'hFFFF;
		end
		32'h0000604C: begin
				q			<=			16'h80E7;
		end
		32'h0000604E: begin
				q			<=			16'h4A80;
		end
		32'h00006050: begin
				q			<=			16'h0863;
		end
		32'h00006052: begin
				q			<=			16'h0005;
		end
		32'h00006054: begin
				q			<=			16'h0593;
		end
		32'h00006056: begin
				q			<=			16'h0009;
		end
		32'h00006058: begin
				q			<=			16'h0513;
		end
		32'h0000605A: begin
				q			<=			16'h0004;
		end
		32'h0000605C: begin
				q			<=			16'hF06F;
		end
		32'h0000605E: begin
				q			<=			16'hFB1F;
		end
		32'h00006060: begin
				q			<=			16'h8513;
		end
		32'h00006062: begin
				q			<=			16'h0004;
		end
		32'h00006064: begin
				q			<=			16'hF097;
		end
		32'h00006066: begin
				q			<=			16'hFFFF;
		end
		32'h00006068: begin
				q			<=			16'h80E7;
		end
		32'h0000606A: begin
				q			<=			16'h6E40;
		end
		32'h0000606C: begin
				q			<=			16'h1A63;
		end
		32'h0000606E: begin
				q			<=			16'h0605;
		end
		32'h00006070: begin
				q			<=			16'h0513;
		end
		32'h00006072: begin
				q			<=			16'h0004;
		end
		32'h00006074: begin
				q			<=			16'hF097;
		end
		32'h00006076: begin
				q			<=			16'hFFFF;
		end
		32'h00006078: begin
				q			<=			16'h80E7;
		end
		32'h0000607A: begin
				q			<=			16'h6D40;
		end
		32'h0000607C: begin
				q			<=			16'h0C63;
		end
		32'h0000607E: begin
				q			<=			16'h0005;
		end
		32'h00006080: begin
				q			<=			16'h9597;
		end
		32'h00006082: begin
				q			<=			16'h0000;
		end
		32'h00006084: begin
				q			<=			16'h8593;
		end
		32'h00006086: begin
				q			<=			16'h22C5;
		end
		32'h00006088: begin
				q			<=			16'h8513;
		end
		32'h0000608A: begin
				q			<=			16'h0004;
		end
		32'h0000608C: begin
				q			<=			16'hF0EF;
		end
		32'h0000608E: begin
				q			<=			16'hDA4F;
		end
		32'h00006090: begin
				q			<=			16'h0263;
		end
		32'h00006092: begin
				q			<=			16'h0605;
		end
		32'h00006094: begin
				q			<=			16'h8513;
		end
		32'h00006096: begin
				q			<=			16'h0004;
		end
		32'h00006098: begin
				q			<=			16'hF097;
		end
		32'h0000609A: begin
				q			<=			16'hFFFF;
		end
		32'h0000609C: begin
				q			<=			16'h80E7;
		end
		32'h0000609E: begin
				q			<=			16'h6B00;
		end
		32'h000060A0: begin
				q			<=			16'h1A63;
		end
		32'h000060A2: begin
				q			<=			16'h0005;
		end
		32'h000060A4: begin
				q			<=			16'h0513;
		end
		32'h000060A6: begin
				q			<=			16'h0004;
		end
		32'h000060A8: begin
				q			<=			16'hF097;
		end
		32'h000060AA: begin
				q			<=			16'hFFFF;
		end
		32'h000060AC: begin
				q			<=			16'h80E7;
		end
		32'h000060AE: begin
				q			<=			16'h6A00;
		end
		32'h000060B0: begin
				q			<=			16'h0E63;
		end
		32'h000060B2: begin
				q			<=			16'h0405;
		end
		32'h000060B4: begin
				q			<=			16'h8513;
		end
		32'h000060B6: begin
				q			<=			16'h0004;
		end
		32'h000060B8: begin
				q			<=			16'hF0EF;
		end
		32'h000060BA: begin
				q			<=			16'hC6CF;
		end
		32'h000060BC: begin
				q			<=			16'h0493;
		end
		32'h000060BE: begin
				q			<=			16'h0005;
		end
		32'h000060C0: begin
				q			<=			16'h0513;
		end
		32'h000060C2: begin
				q			<=			16'h0004;
		end
		32'h000060C4: begin
				q			<=			16'hF0EF;
		end
		32'h000060C6: begin
				q			<=			16'hC60F;
		end
		32'h000060C8: begin
				q			<=			16'h8E63;
		end
		32'h000060CA: begin
				q			<=			16'h02A4;
		end
		32'h000060CC: begin
				q			<=			16'h87B7;
		end
		32'h000060CE: begin
				q			<=			16'hFFFF;
		end
		32'h000060D0: begin
				q			<=			16'h1923;
		end
		32'h000060D2: begin
				q			<=			16'h00F9;
		end
		32'h000060D4: begin
				q			<=			16'h0513;
		end
		32'h000060D6: begin
				q			<=			16'h0009;
		end
		32'h000060D8: begin
				q			<=			16'hF0EF;
		end
		32'h000060DA: begin
				q			<=			16'hEA4F;
		end
		32'h000060DC: begin
				q			<=			16'hF06F;
		end
		32'h000060DE: begin
				q			<=			16'hF35F;
		end
		32'h000060E0: begin
				q			<=			16'h9597;
		end
		32'h000060E2: begin
				q			<=			16'h0000;
		end
		32'h000060E4: begin
				q			<=			16'h8593;
		end
		32'h000060E6: begin
				q			<=			16'h1CC5;
		end
		32'h000060E8: begin
				q			<=			16'h0513;
		end
		32'h000060EA: begin
				q			<=			16'h0004;
		end
		32'h000060EC: begin
				q			<=			16'hF0EF;
		end
		32'h000060EE: begin
				q			<=			16'hD44F;
		end
		32'h000060F0: begin
				q			<=			16'h10E3;
		end
		32'h000060F2: begin
				q			<=			16'hF805;
		end
		32'h000060F4: begin
				q			<=			16'h0513;
		end
		32'h000060F6: begin
				q			<=			16'h0009;
		end
		32'h000060F8: begin
				q			<=			16'h0097;
		end
		32'h000060FA: begin
				q			<=			16'h0000;
		end
		32'h000060FC: begin
				q			<=			16'h80E7;
		end
		32'h000060FE: begin
				q			<=			16'h8F00;
		end
		32'h00006100: begin
				q			<=			16'hF06F;
		end
		32'h00006102: begin
				q			<=			16'hF11F;
		end
		32'h00006104: begin
				q			<=			16'h1923;
		end
		32'h00006106: begin
				q			<=			16'h0009;
		end
		32'h00006108: begin
				q			<=			16'hF06F;
		end
		32'h0000610A: begin
				q			<=			16'hFCDF;
		end
		32'h0000610C: begin
				q			<=			16'h8513;
		end
		32'h0000610E: begin
				q			<=			16'h0004;
		end
		32'h00006110: begin
				q			<=			16'h0593;
		end
		32'h00006112: begin
				q			<=			16'h00C1;
		end
		32'h00006114: begin
				q			<=			16'hF097;
		end
		32'h00006116: begin
				q			<=			16'hFFFF;
		end
		32'h00006118: begin
				q			<=			16'h80E7;
		end
		32'h0000611A: begin
				q			<=			16'h44C0;
		end
		32'h0000611C: begin
				q			<=			16'h0513;
		end
		32'h0000611E: begin
				q			<=			16'h0004;
		end
		32'h00006120: begin
				q			<=			16'h0593;
		end
		32'h00006122: begin
				q			<=			16'h0281;
		end
		32'h00006124: begin
				q			<=			16'hF097;
		end
		32'h00006126: begin
				q			<=			16'hFFFF;
		end
		32'h00006128: begin
				q			<=			16'h80E7;
		end
		32'h0000612A: begin
				q			<=			16'h43C0;
		end
		32'h0000612C: begin
				q			<=			16'h5403;
		end
		32'h0000612E: begin
				q			<=			16'h00E1;
		end
		32'h00006130: begin
				q			<=			16'h5483;
		end
		32'h00006132: begin
				q			<=			16'h02A1;
		end
		32'h00006134: begin
				q			<=			16'h1463;
		end
		32'h00006136: begin
				q			<=			16'h0204;
		end
		32'h00006138: begin
				q			<=			16'h0793;
		end
		32'h0000613A: begin
				q			<=			16'h0000;
		end
		32'h0000613C: begin
				q			<=			16'h0713;
		end
		32'h0000613E: begin
				q			<=			16'h0160;
		end
		32'h00006140: begin
				q			<=			16'h0693;
		end
		32'h00006142: begin
				q			<=			16'h00C1;
		end
		32'h00006144: begin
				q			<=			16'h86B3;
		end
		32'h00006146: begin
				q			<=			16'h00F6;
		end
		32'h00006148: begin
				q			<=			16'hD683;
		end
		32'h0000614A: begin
				q			<=			16'h0026;
		end
		32'h0000614C: begin
				q			<=			16'h8C63;
		end
		32'h0000614E: begin
				q			<=			16'h1006;
		end
		32'h00006150: begin
				q			<=			16'h0513;
		end
		32'h00006152: begin
				q			<=			16'h00C1;
		end
		32'h00006154: begin
				q			<=			16'hF0EF;
		end
		32'h00006156: begin
				q			<=			16'hFB4F;
		end
		32'h00006158: begin
				q			<=			16'h0433;
		end
		32'h0000615A: begin
				q			<=			16'h40A0;
		end
		32'h0000615C: begin
				q			<=			16'h5783;
		end
		32'h0000615E: begin
				q			<=			16'h02A1;
		end
		32'h00006160: begin
				q			<=			16'h8C13;
		end
		32'h00006162: begin
				q			<=			16'h0004;
		end
		32'h00006164: begin
				q			<=			16'h9263;
		end
		32'h00006166: begin
				q			<=			16'h0207;
		end
		32'h00006168: begin
				q			<=			16'h0713;
		end
		32'h0000616A: begin
				q			<=			16'h0160;
		end
		32'h0000616C: begin
				q			<=			16'h0693;
		end
		32'h0000616E: begin
				q			<=			16'h0281;
		end
		32'h00006170: begin
				q			<=			16'h86B3;
		end
		32'h00006172: begin
				q			<=			16'h00F6;
		end
		32'h00006174: begin
				q			<=			16'hD683;
		end
		32'h00006176: begin
				q			<=			16'h0026;
		end
		32'h00006178: begin
				q			<=			16'h8263;
		end
		32'h0000617A: begin
				q			<=			16'h1006;
		end
		32'h0000617C: begin
				q			<=			16'h0513;
		end
		32'h0000617E: begin
				q			<=			16'h0281;
		end
		32'h00006180: begin
				q			<=			16'hF0EF;
		end
		32'h00006182: begin
				q			<=			16'hF88F;
		end
		32'h00006184: begin
				q			<=			16'h8C33;
		end
		32'h00006186: begin
				q			<=			16'h40A4;
		end
		32'h00006188: begin
				q			<=			16'h5783;
		end
		32'h0000618A: begin
				q			<=			16'h0281;
		end
		32'h0000618C: begin
				q			<=			16'h8B93;
		end
		32'h0000618E: begin
				q			<=			16'h0349;
		end
		32'h00006190: begin
				q			<=			16'h8493;
		end
		32'h00006192: begin
				q			<=			16'h0389;
		end
		32'h00006194: begin
				q			<=			16'h9A23;
		end
		32'h00006196: begin
				q			<=			16'h02F9;
		end
		32'h00006198: begin
				q			<=			16'h5783;
		end
		32'h0000619A: begin
				q			<=			16'h02A1;
		end
		32'h0000619C: begin
				q			<=			16'h8A13;
		end
		32'h0000619E: begin
				q			<=			16'h000B;
		end
		32'h000061A0: begin
				q			<=			16'h9B23;
		end
		32'h000061A2: begin
				q			<=			16'h02F9;
		end
		32'h000061A4: begin
				q			<=			16'h8793;
		end
		32'h000061A6: begin
				q			<=			16'h04E9;
		end
		32'h000061A8: begin
				q			<=			16'h9023;
		end
		32'h000061AA: begin
				q			<=			16'h0004;
		end
		32'h000061AC: begin
				q			<=			16'h8493;
		end
		32'h000061AE: begin
				q			<=			16'h0024;
		end
		32'h000061B0: begin
				q			<=			16'h9CE3;
		end
		32'h000061B2: begin
				q			<=			16'hFE97;
		end
		32'h000061B4: begin
				q			<=			16'h0A93;
		end
		32'h000061B6: begin
				q			<=			16'h0000;
		end
		32'h000061B8: begin
				q			<=			16'h0B13;
		end
		32'h000061BA: begin
				q			<=			16'h0000;
		end
		32'h000061BC: begin
				q			<=			16'h0C93;
		end
		32'h000061BE: begin
				q			<=			16'hFEC0;
		end
		32'h000061C0: begin
				q			<=			16'h0793;
		end
		32'h000061C2: begin
				q			<=			16'h00C1;
		end
		32'h000061C4: begin
				q			<=			16'h87B3;
		end
		32'h000061C6: begin
				q			<=			16'h0157;
		end
		32'h000061C8: begin
				q			<=			16'hD503;
		end
		32'h000061CA: begin
				q			<=			16'h0187;
		end
		32'h000061CC: begin
				q			<=			16'h0E63;
		end
		32'h000061CE: begin
				q			<=			16'h0005;
		end
		32'h000061D0: begin
				q			<=			16'h0593;
		end
		32'h000061D2: begin
				q			<=			16'h0281;
		end
		32'h000061D4: begin
				q			<=			16'h0613;
		end
		32'h000061D6: begin
				q			<=			16'h0441;
		end
		32'h000061D8: begin
				q			<=			16'hF0EF;
		end
		32'h000061DA: begin
				q			<=			16'hA7CF;
		end
		32'h000061DC: begin
				q			<=			16'h8593;
		end
		32'h000061DE: begin
				q			<=			16'h000B;
		end
		32'h000061E0: begin
				q			<=			16'h0513;
		end
		32'h000061E2: begin
				q			<=			16'h0441;
		end
		32'h000061E4: begin
				q			<=			16'hF0EF;
		end
		32'h000061E6: begin
				q			<=			16'hA00F;
		end
		32'h000061E8: begin
				q			<=			16'hD783;
		end
		32'h000061EA: begin
				q			<=			16'h04C9;
		end
		32'h000061EC: begin
				q			<=			16'h8513;
		end
		32'h000061EE: begin
				q			<=			16'h000B;
		end
		32'h000061F0: begin
				q			<=			16'h8A93;
		end
		32'h000061F2: begin
				q			<=			16'hFFEA;
		end
		32'h000061F4: begin
				q			<=			16'h6B33;
		end
		32'h000061F6: begin
				q			<=			16'h00FB;
		end
		32'h000061F8: begin
				q			<=			16'hF097;
		end
		32'h000061FA: begin
				q			<=			16'hFFFF;
		end
		32'h000061FC: begin
				q			<=			16'h80E7;
		end
		32'h000061FE: begin
				q			<=			16'h1C40;
		end
		32'h00006200: begin
				q			<=			16'h90E3;
		end
		32'h00006202: begin
				q			<=			16'hFD9A;
		end
		32'h00006204: begin
				q			<=			16'h0793;
		end
		32'h00006206: begin
				q			<=			16'h0281;
		end
		32'h00006208: begin
				q			<=			16'h5703;
		end
		32'h0000620A: begin
				q			<=			16'h000A;
		end
		32'h0000620C: begin
				q			<=			16'h0A13;
		end
		32'h0000620E: begin
				q			<=			16'h002A;
		end
		32'h00006210: begin
				q			<=			16'h8793;
		end
		32'h00006212: begin
				q			<=			16'h0027;
		end
		32'h00006214: begin
				q			<=			16'h9F23;
		end
		32'h00006216: begin
				q			<=			16'hFEE7;
		end
		32'h00006218: begin
				q			<=			16'h18E3;
		end
		32'h0000621A: begin
				q			<=			16'hFE9A;
		end
		32'h0000621C: begin
				q			<=			16'hC6B7;
		end
		32'h0000621E: begin
				q			<=			16'hFFFF;
		end
		32'h00006220: begin
				q			<=			16'h0433;
		end
		32'h00006222: begin
				q			<=			16'h0184;
		end
		32'h00006224: begin
				q			<=			16'h8693;
		end
		32'h00006226: begin
				q			<=			16'h0026;
		end
		32'h00006228: begin
				q			<=			16'h8793;
		end
		32'h0000622A: begin
				q			<=			16'h0009;
		end
		32'h0000622C: begin
				q			<=			16'h0713;
		end
		32'h0000622E: begin
				q			<=			16'h0400;
		end
		32'h00006230: begin
				q			<=			16'h06B3;
		end
		32'h00006232: begin
				q			<=			16'h00D4;
		end
		32'h00006234: begin
				q			<=			16'h0613;
		end
		32'h00006236: begin
				q			<=			16'h0000;
		end
		32'h00006238: begin
				q			<=			16'h0593;
		end
		32'h0000623A: begin
				q			<=			16'h000B;
		end
		32'h0000623C: begin
				q			<=			16'h0513;
		end
		32'h0000623E: begin
				q			<=			16'h0281;
		end
		32'h00006240: begin
				q			<=			16'hF0EF;
		end
		32'h00006242: begin
				q			<=			16'h955F;
		end
		32'h00006244: begin
				q			<=			16'h5703;
		end
		32'h00006246: begin
				q			<=			16'h00C1;
		end
		32'h00006248: begin
				q			<=			16'h5783;
		end
		32'h0000624A: begin
				q			<=			16'h0281;
		end
		32'h0000624C: begin
				q			<=			16'h1E63;
		end
		32'h0000624E: begin
				q			<=			16'h02F7;
		end
		32'h00006250: begin
				q			<=			16'h1423;
		end
		32'h00006252: begin
				q			<=			16'h0201;
		end
		32'h00006254: begin
				q			<=			16'h0593;
		end
		32'h00006256: begin
				q			<=			16'h0009;
		end
		32'h00006258: begin
				q			<=			16'h0513;
		end
		32'h0000625A: begin
				q			<=			16'h0281;
		end
		32'h0000625C: begin
				q			<=			16'hF0EF;
		end
		32'h0000625E: begin
				q			<=			16'hFB4F;
		end
		32'h00006260: begin
				q			<=			16'hF06F;
		end
		32'h00006262: begin
				q			<=			16'hDB1F;
		end
		32'h00006264: begin
				q			<=			16'h8793;
		end
		32'h00006266: begin
				q			<=			16'h0027;
		end
		32'h00006268: begin
				q			<=			16'h9CE3;
		end
		32'h0000626A: begin
				q			<=			16'hECE7;
		end
		32'h0000626C: begin
				q			<=			16'h0513;
		end
		32'h0000626E: begin
				q			<=			16'h0009;
		end
		32'h00006270: begin
				q			<=			16'hF097;
		end
		32'h00006272: begin
				q			<=			16'hFFFF;
		end
		32'h00006274: begin
				q			<=			16'h80E7;
		end
		32'h00006276: begin
				q			<=			16'hF880;
		end
		32'h00006278: begin
				q			<=			16'hF06F;
		end
		32'h0000627A: begin
				q			<=			16'hD99F;
		end
		32'h0000627C: begin
				q			<=			16'h8793;
		end
		32'h0000627E: begin
				q			<=			16'h0027;
		end
		32'h00006280: begin
				q			<=			16'h96E3;
		end
		32'h00006282: begin
				q			<=			16'hEEE7;
		end
		32'h00006284: begin
				q			<=			16'hF06F;
		end
		32'h00006286: begin
				q			<=			16'hFE9F;
		end
		32'h00006288: begin
				q			<=			16'h0793;
		end
		32'h0000628A: begin
				q			<=			16'hFFF0;
		end
		32'h0000628C: begin
				q			<=			16'h1423;
		end
		32'h0000628E: begin
				q			<=			16'h02F1;
		end
		32'h00006290: begin
				q			<=			16'hF06F;
		end
		32'h00006292: begin
				q			<=			16'hFC5F;
		end
		32'h00006294: begin
				q			<=			16'h0113;
		end
		32'h00006296: begin
				q			<=			16'hF701;
		end
		32'h00006298: begin
				q			<=			16'h2423;
		end
		32'h0000629A: begin
				q			<=			16'h0881;
		end
		32'h0000629C: begin
				q			<=			16'h2223;
		end
		32'h0000629E: begin
				q			<=			16'h0891;
		end
		32'h000062A0: begin
				q			<=			16'h2023;
		end
		32'h000062A2: begin
				q			<=			16'h0921;
		end
		32'h000062A4: begin
				q			<=			16'h2A23;
		end
		32'h000062A6: begin
				q			<=			16'h0751;
		end
		32'h000062A8: begin
				q			<=			16'h2623;
		end
		32'h000062AA: begin
				q			<=			16'h0811;
		end
		32'h000062AC: begin
				q			<=			16'h2E23;
		end
		32'h000062AE: begin
				q			<=			16'h0731;
		end
		32'h000062B0: begin
				q			<=			16'h2C23;
		end
		32'h000062B2: begin
				q			<=			16'h0741;
		end
		32'h000062B4: begin
				q			<=			16'h2823;
		end
		32'h000062B6: begin
				q			<=			16'h0761;
		end
		32'h000062B8: begin
				q			<=			16'h2623;
		end
		32'h000062BA: begin
				q			<=			16'h0771;
		end
		32'h000062BC: begin
				q			<=			16'h2423;
		end
		32'h000062BE: begin
				q			<=			16'h0781;
		end
		32'h000062C0: begin
				q			<=			16'h2223;
		end
		32'h000062C2: begin
				q			<=			16'h0791;
		end
		32'h000062C4: begin
				q			<=			16'h2023;
		end
		32'h000062C6: begin
				q			<=			16'h07A1;
		end
		32'h000062C8: begin
				q			<=			16'h0493;
		end
		32'h000062CA: begin
				q			<=			16'h0005;
		end
		32'h000062CC: begin
				q			<=			16'h8413;
		end
		32'h000062CE: begin
				q			<=			16'h0005;
		end
		32'h000062D0: begin
				q			<=			16'h0913;
		end
		32'h000062D2: begin
				q			<=			16'h0006;
		end
		32'h000062D4: begin
				q			<=			16'h8A93;
		end
		32'h000062D6: begin
				q			<=			16'h0006;
		end
		32'h000062D8: begin
				q			<=			16'hF0EF;
		end
		32'h000062DA: begin
				q			<=			16'hA18F;
		end
		32'h000062DC: begin
				q			<=			16'h0663;
		end
		32'h000062DE: begin
				q			<=			16'h0405;
		end
		32'h000062E0: begin
				q			<=			16'h0593;
		end
		32'h000062E2: begin
				q			<=			16'h0009;
		end
		32'h000062E4: begin
				q			<=			16'h8513;
		end
		32'h000062E6: begin
				q			<=			16'h0004;
		end
		32'h000062E8: begin
				q			<=			16'hF097;
		end
		32'h000062EA: begin
				q			<=			16'hFFFF;
		end
		32'h000062EC: begin
				q			<=			16'h80E7;
		end
		32'h000062EE: begin
				q			<=			16'hF240;
		end
		32'h000062F0: begin
				q			<=			16'h2083;
		end
		32'h000062F2: begin
				q			<=			16'h08C1;
		end
		32'h000062F4: begin
				q			<=			16'h2403;
		end
		32'h000062F6: begin
				q			<=			16'h0881;
		end
		32'h000062F8: begin
				q			<=			16'h2483;
		end
		32'h000062FA: begin
				q			<=			16'h0841;
		end
		32'h000062FC: begin
				q			<=			16'h2903;
		end
		32'h000062FE: begin
				q			<=			16'h0801;
		end
		32'h00006300: begin
				q			<=			16'h2983;
		end
		32'h00006302: begin
				q			<=			16'h07C1;
		end
		32'h00006304: begin
				q			<=			16'h2A03;
		end
		32'h00006306: begin
				q			<=			16'h0781;
		end
		32'h00006308: begin
				q			<=			16'h2A83;
		end
		32'h0000630A: begin
				q			<=			16'h0741;
		end
		32'h0000630C: begin
				q			<=			16'h2B03;
		end
		32'h0000630E: begin
				q			<=			16'h0701;
		end
		32'h00006310: begin
				q			<=			16'h2B83;
		end
		32'h00006312: begin
				q			<=			16'h06C1;
		end
		32'h00006314: begin
				q			<=			16'h2C03;
		end
		32'h00006316: begin
				q			<=			16'h0681;
		end
		32'h00006318: begin
				q			<=			16'h2C83;
		end
		32'h0000631A: begin
				q			<=			16'h0641;
		end
		32'h0000631C: begin
				q			<=			16'h2D03;
		end
		32'h0000631E: begin
				q			<=			16'h0601;
		end
		32'h00006320: begin
				q			<=			16'h0113;
		end
		32'h00006322: begin
				q			<=			16'h0901;
		end
		32'h00006324: begin
				q			<=			16'h8067;
		end
		32'h00006326: begin
				q			<=			16'h0000;
		end
		32'h00006328: begin
				q			<=			16'h0513;
		end
		32'h0000632A: begin
				q			<=			16'h0004;
		end
		32'h0000632C: begin
				q			<=			16'hF0EF;
		end
		32'h0000632E: begin
				q			<=			16'h9C4F;
		end
		32'h00006330: begin
				q			<=			16'h0863;
		end
		32'h00006332: begin
				q			<=			16'h0005;
		end
		32'h00006334: begin
				q			<=			16'h0593;
		end
		32'h00006336: begin
				q			<=			16'h0009;
		end
		32'h00006338: begin
				q			<=			16'h0513;
		end
		32'h0000633A: begin
				q			<=			16'h0004;
		end
		32'h0000633C: begin
				q			<=			16'hF06F;
		end
		32'h0000633E: begin
				q			<=			16'hFADF;
		end
		32'h00006340: begin
				q			<=			16'h9597;
		end
		32'h00006342: begin
				q			<=			16'h0000;
		end
		32'h00006344: begin
				q			<=			16'h8593;
		end
		32'h00006346: begin
				q			<=			16'hF6C5;
		end
		32'h00006348: begin
				q			<=			16'h8513;
		end
		32'h0000634A: begin
				q			<=			16'h0004;
		end
		32'h0000634C: begin
				q			<=			16'hF097;
		end
		32'h0000634E: begin
				q			<=			16'hFFFF;
		end
		32'h00006350: begin
				q			<=			16'h80E7;
		end
		32'h00006352: begin
				q			<=			16'h2E40;
		end
		32'h00006354: begin
				q			<=			16'h0463;
		end
		32'h00006356: begin
				q			<=			16'h2005;
		end
		32'h00006358: begin
				q			<=			16'h8513;
		end
		32'h0000635A: begin
				q			<=			16'h0004;
		end
		32'h0000635C: begin
				q			<=			16'hF0EF;
		end
		32'h0000635E: begin
				q			<=			16'hBECF;
		end
		32'h00006360: begin
				q			<=			16'h0993;
		end
		32'h00006362: begin
				q			<=			16'h0005;
		end
		32'h00006364: begin
				q			<=			16'h0513;
		end
		32'h00006366: begin
				q			<=			16'h0004;
		end
		32'h00006368: begin
				q			<=			16'hF0EF;
		end
		32'h0000636A: begin
				q			<=			16'hBE0F;
		end
		32'h0000636C: begin
				q			<=			16'h9A63;
		end
		32'h0000636E: begin
				q			<=			16'h2009;
		end
		32'h00006370: begin
				q			<=			16'h1063;
		end
		32'h00006372: begin
				q			<=			16'h2205;
		end
		32'h00006374: begin
				q			<=			16'h8513;
		end
		32'h00006376: begin
				q			<=			16'h0004;
		end
		32'h00006378: begin
				q			<=			16'h0593;
		end
		32'h0000637A: begin
				q			<=			16'h00C1;
		end
		32'h0000637C: begin
				q			<=			16'hF0EF;
		end
		32'h0000637E: begin
				q			<=			16'h9E4F;
		end
		32'h00006380: begin
				q			<=			16'h0513;
		end
		32'h00006382: begin
				q			<=			16'h0004;
		end
		32'h00006384: begin
				q			<=			16'h0593;
		end
		32'h00006386: begin
				q			<=			16'h0281;
		end
		32'h00006388: begin
				q			<=			16'hF0EF;
		end
		32'h0000638A: begin
				q			<=			16'h9D8F;
		end
		32'h0000638C: begin
				q			<=			16'h5483;
		end
		32'h0000638E: begin
				q			<=			16'h02A1;
		end
		32'h00006390: begin
				q			<=			16'h5403;
		end
		32'h00006392: begin
				q			<=			16'h00E1;
		end
		32'h00006394: begin
				q			<=			16'h9663;
		end
		32'h00006396: begin
				q			<=			16'h0204;
		end
		32'h00006398: begin
				q			<=			16'h0793;
		end
		32'h0000639A: begin
				q			<=			16'h0000;
		end
		32'h0000639C: begin
				q			<=			16'h0713;
		end
		32'h0000639E: begin
				q			<=			16'h0160;
		end
		32'h000063A0: begin
				q			<=			16'h0693;
		end
		32'h000063A2: begin
				q			<=			16'h0281;
		end
		32'h000063A4: begin
				q			<=			16'h86B3;
		end
		32'h000063A6: begin
				q			<=			16'h00F6;
		end
		32'h000063A8: begin
				q			<=			16'hD683;
		end
		32'h000063AA: begin
				q			<=			16'h0026;
		end
		32'h000063AC: begin
				q			<=			16'h8E63;
		end
		32'h000063AE: begin
				q			<=			16'h2006;
		end
		32'h000063B0: begin
				q			<=			16'h0513;
		end
		32'h000063B2: begin
				q			<=			16'h0281;
		end
		32'h000063B4: begin
				q			<=			16'hF097;
		end
		32'h000063B6: begin
				q			<=			16'hFFFF;
		end
		32'h000063B8: begin
				q			<=			16'h80E7;
		end
		32'h000063BA: begin
				q			<=			16'h5540;
		end
		32'h000063BC: begin
				q			<=			16'h04B3;
		end
		32'h000063BE: begin
				q			<=			16'h40A0;
		end
		32'h000063C0: begin
				q			<=			16'h5783;
		end
		32'h000063C2: begin
				q			<=			16'h00E1;
		end
		32'h000063C4: begin
				q			<=			16'h0B93;
		end
		32'h000063C6: begin
				q			<=			16'h0004;
		end
		32'h000063C8: begin
				q			<=			16'h9463;
		end
		32'h000063CA: begin
				q			<=			16'h0207;
		end
		32'h000063CC: begin
				q			<=			16'h0713;
		end
		32'h000063CE: begin
				q			<=			16'h0160;
		end
		32'h000063D0: begin
				q			<=			16'h0693;
		end
		32'h000063D2: begin
				q			<=			16'h00C1;
		end
		32'h000063D4: begin
				q			<=			16'h86B3;
		end
		32'h000063D6: begin
				q			<=			16'h00F6;
		end
		32'h000063D8: begin
				q			<=			16'hD683;
		end
		32'h000063DA: begin
				q			<=			16'h0026;
		end
		32'h000063DC: begin
				q			<=			16'h8C63;
		end
		32'h000063DE: begin
				q			<=			16'h1E06;
		end
		32'h000063E0: begin
				q			<=			16'h0513;
		end
		32'h000063E2: begin
				q			<=			16'h00C1;
		end
		32'h000063E4: begin
				q			<=			16'hF097;
		end
		32'h000063E6: begin
				q			<=			16'hFFFF;
		end
		32'h000063E8: begin
				q			<=			16'h80E7;
		end
		32'h000063EA: begin
				q			<=			16'h5240;
		end
		32'h000063EC: begin
				q			<=			16'h0BB3;
		end
		32'h000063EE: begin
				q			<=			16'h40A4;
		end
		32'h000063F0: begin
				q			<=			16'h5783;
		end
		32'h000063F2: begin
				q			<=			16'h0281;
		end
		32'h000063F4: begin
				q			<=			16'h5703;
		end
		32'h000063F6: begin
				q			<=			16'h02A1;
		end
		32'h000063F8: begin
				q			<=			16'h8993;
		end
		32'h000063FA: begin
				q			<=			16'h034A;
		end
		32'h000063FC: begin
				q			<=			16'h9A23;
		end
		32'h000063FE: begin
				q			<=			16'h02FA;
		end
		32'h00006400: begin
				q			<=			16'h8793;
		end
		32'h00006402: begin
				q			<=			16'h038A;
		end
		32'h00006404: begin
				q			<=			16'h9B23;
		end
		32'h00006406: begin
				q			<=			16'h02EA;
		end
		32'h00006408: begin
				q			<=			16'h8A13;
		end
		32'h0000640A: begin
				q			<=			16'h0007;
		end
		32'h0000640C: begin
				q			<=			16'h8713;
		end
		32'h0000640E: begin
				q			<=			16'h04EA;
		end
		32'h00006410: begin
				q			<=			16'h8793;
		end
		32'h00006412: begin
				q			<=			16'h0027;
		end
		32'h00006414: begin
				q			<=			16'h9F23;
		end
		32'h00006416: begin
				q			<=			16'hFE07;
		end
		32'h00006418: begin
				q			<=			16'h9CE3;
		end
		32'h0000641A: begin
				q			<=			16'hFEE7;
		end
		32'h0000641C: begin
				q			<=			16'h0513;
		end
		32'h0000641E: begin
				q			<=			16'h0281;
		end
		32'h00006420: begin
				q			<=			16'hF097;
		end
		32'h00006422: begin
				q			<=			16'hFFFF;
		end
		32'h00006424: begin
				q			<=			16'h80E7;
		end
		32'h00006426: begin
				q			<=			16'hE7C0;
		end
		32'h00006428: begin
				q			<=			16'h5C03;
		end
		32'h0000642A: begin
				q			<=			16'h0121;
		end
		32'h0000642C: begin
				q			<=			16'h0B37;
		end
		32'h0000642E: begin
				q			<=			16'h0001;
		end
		32'h00006430: begin
				q			<=			16'h0B13;
		end
		32'h00006432: begin
				q			<=			16'hFFFB;
		end
		32'h00006434: begin
				q			<=			16'h0D33;
		end
		32'h00006436: begin
				q			<=			16'h036C;
		end
		32'h00006438: begin
				q			<=			16'h8C93;
		end
		32'h0000643A: begin
				q			<=			16'h01A9;
		end
		32'h0000643C: begin
				q			<=			16'h5783;
		end
		32'h0000643E: begin
				q			<=			16'h02C1;
		end
		32'h00006440: begin
				q			<=			16'h5403;
		end
		32'h00006442: begin
				q			<=			16'h02E1;
		end
		32'h00006444: begin
				q			<=			16'h9793;
		end
		32'h00006446: begin
				q			<=			16'h0107;
		end
		32'h00006448: begin
				q			<=			16'h87B3;
		end
		32'h0000644A: begin
				q			<=			16'h0087;
		end
		32'h0000644C: begin
				q			<=			16'h0413;
		end
		32'h0000644E: begin
				q			<=			16'h000B;
		end
		32'h00006450: begin
				q			<=			16'h6863;
		end
		32'h00006452: begin
				q			<=			16'h00FD;
		end
		32'h00006454: begin
				q			<=			16'hD433;
		end
		32'h00006456: begin
				q			<=			16'h0387;
		end
		32'h00006458: begin
				q			<=			16'h1413;
		end
		32'h0000645A: begin
				q			<=			16'h0104;
		end
		32'h0000645C: begin
				q			<=			16'h5413;
		end
		32'h0000645E: begin
				q			<=			16'h0104;
		end
		32'h00006460: begin
				q			<=			16'h0593;
		end
		32'h00006462: begin
				q			<=			16'h00C1;
		end
		32'h00006464: begin
				q			<=			16'h0513;
		end
		32'h00006466: begin
				q			<=			16'h0004;
		end
		32'h00006468: begin
				q			<=			16'h0613;
		end
		32'h0000646A: begin
				q			<=			16'h0441;
		end
		32'h0000646C: begin
				q			<=			16'hF097;
		end
		32'h0000646E: begin
				q			<=			16'hFFFF;
		end
		32'h00006470: begin
				q			<=			16'h80E7;
		end
		32'h00006472: begin
				q			<=			16'hFE80;
		end
		32'h00006474: begin
				q			<=			16'h0593;
		end
		32'h00006476: begin
				q			<=			16'h0281;
		end
		32'h00006478: begin
				q			<=			16'h0513;
		end
		32'h0000647A: begin
				q			<=			16'h0441;
		end
		32'h0000647C: begin
				q			<=			16'hE0EF;
		end
		32'h0000647E: begin
				q			<=			16'hDE5F;
		end
		32'h00006480: begin
				q			<=			16'h5663;
		end
		32'h00006482: begin
				q			<=			16'h02A0;
		end
		32'h00006484: begin
				q			<=			16'h0593;
		end
		32'h00006486: begin
				q			<=			16'h0441;
		end
		32'h00006488: begin
				q			<=			16'h0513;
		end
		32'h0000648A: begin
				q			<=			16'h00C1;
		end
		32'h0000648C: begin
				q			<=			16'hE0EF;
		end
		32'h0000648E: begin
				q			<=			16'hF91F;
		end
		32'h00006490: begin
				q			<=			16'h0593;
		end
		32'h00006492: begin
				q			<=			16'h0281;
		end
		32'h00006494: begin
				q			<=			16'h0513;
		end
		32'h00006496: begin
				q			<=			16'h0441;
		end
		32'h00006498: begin
				q			<=			16'hE0EF;
		end
		32'h0000649A: begin
				q			<=			16'hDC9F;
		end
		32'h0000649C: begin
				q			<=			16'h4A63;
		end
		32'h0000649E: begin
				q			<=			16'h14A0;
		end
		32'h000064A0: begin
				q			<=			16'h0413;
		end
		32'h000064A2: begin
				q			<=			16'hFFF4;
		end
		32'h000064A4: begin
				q			<=			16'h1413;
		end
		32'h000064A6: begin
				q			<=			16'h0104;
		end
		32'h000064A8: begin
				q			<=			16'h5413;
		end
		32'h000064AA: begin
				q			<=			16'h0104;
		end
		32'h000064AC: begin
				q			<=			16'h0593;
		end
		32'h000064AE: begin
				q			<=			16'h0281;
		end
		32'h000064B0: begin
				q			<=			16'h0513;
		end
		32'h000064B2: begin
				q			<=			16'h0441;
		end
		32'h000064B4: begin
				q			<=			16'hE0EF;
		end
		32'h000064B6: begin
				q			<=			16'hF69F;
		end
		32'h000064B8: begin
				q			<=			16'h0513;
		end
		32'h000064BA: begin
				q			<=			16'h0281;
		end
		32'h000064BC: begin
				q			<=			16'h1023;
		end
		32'h000064BE: begin
				q			<=			16'h008A;
		end
		32'h000064C0: begin
				q			<=			16'h0A13;
		end
		32'h000064C2: begin
				q			<=			16'h002A;
		end
		32'h000064C4: begin
				q			<=			16'hF097;
		end
		32'h000064C6: begin
				q			<=			16'hFFFF;
		end
		32'h000064C8: begin
				q			<=			16'h80E7;
		end
		32'h000064CA: begin
				q			<=			16'hED80;
		end
		32'h000064CC: begin
				q			<=			16'h18E3;
		end
		32'h000064CE: begin
				q			<=			16'hF79A;
		end
		32'h000064D0: begin
				q			<=			16'h0793;
		end
		32'h000064D2: begin
				q			<=			16'h0000;
		end
		32'h000064D4: begin
				q			<=			16'h0593;
		end
		32'h000064D6: begin
				q			<=			16'h0000;
		end
		32'h000064D8: begin
				q			<=			16'h0713;
		end
		32'h000064DA: begin
				q			<=			16'h0160;
		end
		32'h000064DC: begin
				q			<=			16'h0693;
		end
		32'h000064DE: begin
				q			<=			16'h0281;
		end
		32'h000064E0: begin
				q			<=			16'h86B3;
		end
		32'h000064E2: begin
				q			<=			16'h00F6;
		end
		32'h000064E4: begin
				q			<=			16'hD683;
		end
		32'h000064E6: begin
				q			<=			16'h0046;
		end
		32'h000064E8: begin
				q			<=			16'h8793;
		end
		32'h000064EA: begin
				q			<=			16'h0027;
		end
		32'h000064EC: begin
				q			<=			16'hE5B3;
		end
		32'h000064EE: begin
				q			<=			16'h00D5;
		end
		32'h000064F0: begin
				q			<=			16'h96E3;
		end
		32'h000064F2: begin
				q			<=			16'hFEE7;
		end
		32'h000064F4: begin
				q			<=			16'h35B3;
		end
		32'h000064F6: begin
				q			<=			16'h00B0;
		end
		32'h000064F8: begin
				q			<=			16'h0793;
		end
		32'h000064FA: begin
				q			<=			16'h0281;
		end
		32'h000064FC: begin
				q			<=			16'hD703;
		end
		32'h000064FE: begin
				q			<=			16'h0009;
		end
		32'h00006500: begin
				q			<=			16'h8993;
		end
		32'h00006502: begin
				q			<=			16'h0029;
		end
		32'h00006504: begin
				q			<=			16'h8793;
		end
		32'h00006506: begin
				q			<=			16'h0027;
		end
		32'h00006508: begin
				q			<=			16'h9F23;
		end
		32'h0000650A: begin
				q			<=			16'hFEE7;
		end
		32'h0000650C: begin
				q			<=			16'h18E3;
		end
		32'h0000650E: begin
				q			<=			16'hFF3A;
		end
		32'h00006510: begin
				q			<=			16'h46B7;
		end
		32'h00006512: begin
				q			<=			16'h0000;
		end
		32'h00006514: begin
				q			<=			16'h84B3;
		end
		32'h00006516: begin
				q			<=			16'h4174;
		end
		32'h00006518: begin
				q			<=			16'h8693;
		end
		32'h0000651A: begin
				q			<=			16'hFFF6;
		end
		32'h0000651C: begin
				q			<=			16'h8793;
		end
		32'h0000651E: begin
				q			<=			16'h000A;
		end
		32'h00006520: begin
				q			<=			16'h0713;
		end
		32'h00006522: begin
				q			<=			16'h0400;
		end
		32'h00006524: begin
				q			<=			16'h86B3;
		end
		32'h00006526: begin
				q			<=			16'h00D4;
		end
		32'h00006528: begin
				q			<=			16'h0613;
		end
		32'h0000652A: begin
				q			<=			16'h0000;
		end
		32'h0000652C: begin
				q			<=			16'h0513;
		end
		32'h0000652E: begin
				q			<=			16'h0281;
		end
		32'h00006530: begin
				q			<=			16'hF097;
		end
		32'h00006532: begin
				q			<=			16'hFFFF;
		end
		32'h00006534: begin
				q			<=			16'h80E7;
		end
		32'h00006536: begin
				q			<=			16'h6640;
		end
		32'h00006538: begin
				q			<=			16'h5703;
		end
		32'h0000653A: begin
				q			<=			16'h00C1;
		end
		32'h0000653C: begin
				q			<=			16'h5783;
		end
		32'h0000653E: begin
				q			<=			16'h0281;
		end
		32'h00006540: begin
				q			<=			16'h1663;
		end
		32'h00006542: begin
				q			<=			16'h0CF7;
		end
		32'h00006544: begin
				q			<=			16'h1423;
		end
		32'h00006546: begin
				q			<=			16'h0201;
		end
		32'h00006548: begin
				q			<=			16'h0593;
		end
		32'h0000654A: begin
				q			<=			16'h0009;
		end
		32'h0000654C: begin
				q			<=			16'h0513;
		end
		32'h0000654E: begin
				q			<=			16'h0281;
		end
		32'h00006550: begin
				q			<=			16'hF097;
		end
		32'h00006552: begin
				q			<=			16'hFFFF;
		end
		32'h00006554: begin
				q			<=			16'h80E7;
		end
		32'h00006556: begin
				q			<=			16'h4C00;
		end
		32'h00006558: begin
				q			<=			16'hF06F;
		end
		32'h0000655A: begin
				q			<=			16'hD99F;
		end
		32'h0000655C: begin
				q			<=			16'h9597;
		end
		32'h0000655E: begin
				q			<=			16'h0000;
		end
		32'h00006560: begin
				q			<=			16'h8593;
		end
		32'h00006562: begin
				q			<=			16'hD505;
		end
		32'h00006564: begin
				q			<=			16'h0513;
		end
		32'h00006566: begin
				q			<=			16'h0004;
		end
		32'h00006568: begin
				q			<=			16'hF097;
		end
		32'h0000656A: begin
				q			<=			16'hFFFF;
		end
		32'h0000656C: begin
				q			<=			16'h80E7;
		end
		32'h0000656E: begin
				q			<=			16'h0C80;
		end
		32'h00006570: begin
				q			<=			16'h14E3;
		end
		32'h00006572: begin
				q			<=			16'hDE05;
		end
		32'h00006574: begin
				q			<=			16'h0513;
		end
		32'h00006576: begin
				q			<=			16'h0009;
		end
		32'h00006578: begin
				q			<=			16'hF0EF;
		end
		32'h0000657A: begin
				q			<=			16'hC70F;
		end
		32'h0000657C: begin
				q			<=			16'hF06F;
		end
		32'h0000657E: begin
				q			<=			16'hD75F;
		end
		32'h00006580: begin
				q			<=			16'h1AE3;
		end
		32'h00006582: begin
				q			<=			16'hFE05;
		end
		32'h00006584: begin
				q			<=			16'h0513;
		end
		32'h00006586: begin
				q			<=			16'h0009;
		end
		32'h00006588: begin
				q			<=			16'hE0EF;
		end
		32'h0000658A: begin
				q			<=			16'hC71F;
		end
		32'h0000658C: begin
				q			<=			16'hF06F;
		end
		32'h0000658E: begin
				q			<=			16'hD65F;
		end
		32'h00006590: begin
				q			<=			16'h8513;
		end
		32'h00006592: begin
				q			<=			16'h0004;
		end
		32'h00006594: begin
				q			<=			16'hF097;
		end
		32'h00006596: begin
				q			<=			16'hFFFF;
		end
		32'h00006598: begin
				q			<=			16'h80E7;
		end
		32'h0000659A: begin
				q			<=			16'hF900;
		end
		32'h0000659C: begin
				q			<=			16'h0493;
		end
		32'h0000659E: begin
				q			<=			16'h0005;
		end
		32'h000065A0: begin
				q			<=			16'h0513;
		end
		32'h000065A2: begin
				q			<=			16'h0004;
		end
		32'h000065A4: begin
				q			<=			16'hF097;
		end
		32'h000065A6: begin
				q			<=			16'hFFFF;
		end
		32'h000065A8: begin
				q			<=			16'h80E7;
		end
		32'h000065AA: begin
				q			<=			16'hF800;
		end
		32'h000065AC: begin
				q			<=			16'h8E63;
		end
		32'h000065AE: begin
				q			<=			16'h02A4;
		end
		32'h000065B0: begin
				q			<=			16'h87B7;
		end
		32'h000065B2: begin
				q			<=			16'hFFFF;
		end
		32'h000065B4: begin
				q			<=			16'h1923;
		end
		32'h000065B6: begin
				q			<=			16'h00F9;
		end
		32'h000065B8: begin
				q			<=			16'h0513;
		end
		32'h000065BA: begin
				q			<=			16'h0009;
		end
		32'h000065BC: begin
				q			<=			16'hF097;
		end
		32'h000065BE: begin
				q			<=			16'hFFFF;
		end
		32'h000065C0: begin
				q			<=			16'h80E7;
		end
		32'h000065C2: begin
				q			<=			16'h1C00;
		end
		32'h000065C4: begin
				q			<=			16'hF06F;
		end
		32'h000065C6: begin
				q			<=			16'hD2DF;
		end
		32'h000065C8: begin
				q			<=			16'h8793;
		end
		32'h000065CA: begin
				q			<=			16'h0027;
		end
		32'h000065CC: begin
				q			<=			16'h9AE3;
		end
		32'h000065CE: begin
				q			<=			16'hDCE7;
		end
		32'h000065D0: begin
				q			<=			16'hF06F;
		end
		32'h000065D2: begin
				q			<=			16'hFB5F;
		end
		32'h000065D4: begin
				q			<=			16'h8793;
		end
		32'h000065D6: begin
				q			<=			16'h0027;
		end
		32'h000065D8: begin
				q			<=			16'h9CE3;
		end
		32'h000065DA: begin
				q			<=			16'hDEE7;
		end
		32'h000065DC: begin
				q			<=			16'h5703;
		end
		32'h000065DE: begin
				q			<=			16'h00C1;
		end
		32'h000065E0: begin
				q			<=			16'h5783;
		end
		32'h000065E2: begin
				q			<=			16'h0281;
		end
		32'h000065E4: begin
				q			<=			16'h16E3;
		end
		32'h000065E6: begin
				q			<=			16'hFCF7;
		end
		32'h000065E8: begin
				q			<=			16'h1923;
		end
		32'h000065EA: begin
				q			<=			16'h0009;
		end
		32'h000065EC: begin
				q			<=			16'hF06F;
		end
		32'h000065EE: begin
				q			<=			16'hFCDF;
		end
		32'h000065F0: begin
				q			<=			16'h0413;
		end
		32'h000065F2: begin
				q			<=			16'hFFE4;
		end
		32'h000065F4: begin
				q			<=			16'h1413;
		end
		32'h000065F6: begin
				q			<=			16'h0104;
		end
		32'h000065F8: begin
				q			<=			16'h0593;
		end
		32'h000065FA: begin
				q			<=			16'h0441;
		end
		32'h000065FC: begin
				q			<=			16'h0513;
		end
		32'h000065FE: begin
				q			<=			16'h00C1;
		end
		32'h00006600: begin
				q			<=			16'h5413;
		end
		32'h00006602: begin
				q			<=			16'h0104;
		end
		32'h00006604: begin
				q			<=			16'hE0EF;
		end
		32'h00006606: begin
				q			<=			16'hE19F;
		end
		32'h00006608: begin
				q			<=			16'hF06F;
		end
		32'h0000660A: begin
				q			<=			16'hEA5F;
		end
		32'h0000660C: begin
				q			<=			16'h0793;
		end
		32'h0000660E: begin
				q			<=			16'hFFF0;
		end
		32'h00006610: begin
				q			<=			16'h1423;
		end
		32'h00006612: begin
				q			<=			16'h02F1;
		end
		32'h00006614: begin
				q			<=			16'hF06F;
		end
		32'h00006616: begin
				q			<=			16'hF35F;
		end
		32'h00006618: begin
				q			<=			16'hAE03;
		end
		32'h0000661A: begin
				q			<=			16'h0005;
		end
		32'h0000661C: begin
				q			<=			16'hA303;
		end
		32'h0000661E: begin
				q			<=			16'h0045;
		end
		32'h00006620: begin
				q			<=			16'hA883;
		end
		32'h00006622: begin
				q			<=			16'h0085;
		end
		32'h00006624: begin
				q			<=			16'hA583;
		end
		32'h00006626: begin
				q			<=			16'h00C5;
		end
		32'h00006628: begin
				q			<=			16'h0113;
		end
		32'h0000662A: begin
				q			<=			16'hE201;
		end
		32'h0000662C: begin
				q			<=			16'h2C23;
		end
		32'h0000662E: begin
				q			<=			16'h1C81;
		end
		32'h00006630: begin
				q			<=			16'h2623;
		end
		32'h00006632: begin
				q			<=			16'h02B1;
		end
		32'h00006634: begin
				q			<=			16'h8413;
		end
		32'h00006636: begin
				q			<=			16'h0007;
		end
		32'h00006638: begin
				q			<=			16'h2583;
		end
		32'h0000663A: begin
				q			<=			16'h0405;
		end
		32'h0000663C: begin
				q			<=			16'h0793;
		end
		32'h0000663E: begin
				q			<=			16'hFFF0;
		end
		32'h00006640: begin
				q			<=			16'h2823;
		end
		32'h00006642: begin
				q			<=			16'h14F1;
		end
		32'h00006644: begin
				q			<=			16'h0793;
		end
		32'h00006646: begin
				q			<=			16'h0900;
		end
		32'h00006648: begin
				q			<=			16'h2823;
		end
		32'h0000664A: begin
				q			<=			16'h1D21;
		end
		32'h0000664C: begin
				q			<=			16'h2623;
		end
		32'h0000664E: begin
				q			<=			16'h1D31;
		end
		32'h00006650: begin
				q			<=			16'h2423;
		end
		32'h00006652: begin
				q			<=			16'h1D41;
		end
		32'h00006654: begin
				q			<=			16'h2E23;
		end
		32'h00006656: begin
				q			<=			16'h1B71;
		end
		32'h00006658: begin
				q			<=			16'h2E23;
		end
		32'h0000665A: begin
				q			<=			16'h1C11;
		end
		32'h0000665C: begin
				q			<=			16'h2A23;
		end
		32'h0000665E: begin
				q			<=			16'h1C91;
		end
		32'h00006660: begin
				q			<=			16'h2223;
		end
		32'h00006662: begin
				q			<=			16'h1D51;
		end
		32'h00006664: begin
				q			<=			16'h2023;
		end
		32'h00006666: begin
				q			<=			16'h1D61;
		end
		32'h00006668: begin
				q			<=			16'h2C23;
		end
		32'h0000666A: begin
				q			<=			16'h1B81;
		end
		32'h0000666C: begin
				q			<=			16'h2A23;
		end
		32'h0000666E: begin
				q			<=			16'h1B91;
		end
		32'h00006670: begin
				q			<=			16'h2823;
		end
		32'h00006672: begin
				q			<=			16'h1BA1;
		end
		32'h00006674: begin
				q			<=			16'h2623;
		end
		32'h00006676: begin
				q			<=			16'h1BB1;
		end
		32'h00006678: begin
				q			<=			16'h2623;
		end
		32'h0000667A: begin
				q			<=			16'h0101;
		end
		32'h0000667C: begin
				q			<=			16'h2023;
		end
		32'h0000667E: begin
				q			<=			16'h03C1;
		end
		32'h00006680: begin
				q			<=			16'h2223;
		end
		32'h00006682: begin
				q			<=			16'h0261;
		end
		32'h00006684: begin
				q			<=			16'h2423;
		end
		32'h00006686: begin
				q			<=			16'h0311;
		end
		32'h00006688: begin
				q			<=			16'h2A23;
		end
		32'h0000668A: begin
				q			<=			16'h14F1;
		end
		32'h0000668C: begin
				q			<=			16'h0913;
		end
		32'h0000668E: begin
				q			<=			16'h0005;
		end
		32'h00006690: begin
				q			<=			16'h0A13;
		end
		32'h00006692: begin
				q			<=			16'h0006;
		end
		32'h00006694: begin
				q			<=			16'h8993;
		end
		32'h00006696: begin
				q			<=			16'h0006;
		end
		32'h00006698: begin
				q			<=			16'h0B93;
		end
		32'h0000669A: begin
				q			<=			16'h0007;
		end
		32'h0000669C: begin
				q			<=			16'h8063;
		end
		32'h0000669E: begin
				q			<=			16'h0205;
		end
		32'h000066A0: begin
				q			<=			16'h2783;
		end
		32'h000066A2: begin
				q			<=			16'h0445;
		end
		32'h000066A4: begin
				q			<=			16'h0713;
		end
		32'h000066A6: begin
				q			<=			16'h0010;
		end
		32'h000066A8: begin
				q			<=			16'h1733;
		end
		32'h000066AA: begin
				q			<=			16'h00F7;
		end
		32'h000066AC: begin
				q			<=			16'hA223;
		end
		32'h000066AE: begin
				q			<=			16'h00F5;
		end
		32'h000066B0: begin
				q			<=			16'hA423;
		end
		32'h000066B2: begin
				q			<=			16'h00E5;
		end
		32'h000066B4: begin
				q			<=			16'h10EF;
		end
		32'h000066B6: begin
				q			<=			16'h4800;
		end
		32'h000066B8: begin
				q			<=			16'h2023;
		end
		32'h000066BA: begin
				q			<=			16'h0409;
		end
		32'h000066BC: begin
				q			<=			16'h0513;
		end
		32'h000066BE: begin
				q			<=			16'h0201;
		end
		32'h000066C0: begin
				q			<=			16'h0593;
		end
		32'h000066C2: begin
				q			<=			16'h0501;
		end
		32'h000066C4: begin
				q			<=			16'hF097;
		end
		32'h000066C6: begin
				q			<=			16'hFFFF;
		end
		32'h000066C8: begin
				q			<=			16'h80E7;
		end
		32'h000066CA: begin
				q			<=			16'h3C00;
		end
		32'h000066CC: begin
				q			<=			16'h0513;
		end
		32'h000066CE: begin
				q			<=			16'h0501;
		end
		32'h000066D0: begin
				q			<=			16'hE0EF;
		end
		32'h000066D2: begin
				q			<=			16'hE55F;
		end
		32'h000066D4: begin
				q			<=			16'h0663;
		end
		32'h000066D6: begin
				q			<=			16'h1A05;
		end
		32'h000066D8: begin
				q			<=			16'h0793;
		end
		32'h000066DA: begin
				q			<=			16'h0010;
		end
		32'h000066DC: begin
				q			<=			16'h2023;
		end
		32'h000066DE: begin
				q			<=			16'h00F4;
		end
		32'h000066E0: begin
				q			<=			16'h0793;
		end
		32'h000066E2: begin
				q			<=			16'h0030;
		end
		32'h000066E4: begin
				q			<=			16'h0263;
		end
		32'h000066E6: begin
				q			<=			16'h1AFA;
		end
		32'h000066E8: begin
				q			<=			16'h0493;
		end
		32'h000066EA: begin
				q			<=			16'h0140;
		end
		32'h000066EC: begin
				q			<=			16'h0A63;
		end
		32'h000066EE: begin
				q			<=			16'h000A;
		end
		32'h000066F0: begin
				q			<=			16'h8493;
		end
		32'h000066F2: begin
				q			<=			16'hFFF9;
		end
		32'h000066F4: begin
				q			<=			16'h0793;
		end
		32'h000066F6: begin
				q			<=			16'h02A0;
		end
		32'h000066F8: begin
				q			<=			16'hD463;
		end
		32'h000066FA: begin
				q			<=			16'h0097;
		end
		32'h000066FC: begin
				q			<=			16'h0493;
		end
		32'h000066FE: begin
				q			<=			16'h02A0;
		end
		32'h00006700: begin
				q			<=			16'h2783;
		end
		32'h00006702: begin
				q			<=			16'h1541;
		end
		32'h00006704: begin
				q			<=			16'h0513;
		end
		32'h00006706: begin
				q			<=			16'h0501;
		end
		32'h00006708: begin
				q			<=			16'h2823;
		end
		32'h0000670A: begin
				q			<=			16'h00F1;
		end
		32'h0000670C: begin
				q			<=			16'hF097;
		end
		32'h0000670E: begin
				q			<=			16'hFFFF;
		end
		32'h00006710: begin
				q			<=			16'h80E7;
		end
		32'h00006712: begin
				q			<=			16'hDE40;
		end
		32'h00006714: begin
				q			<=			16'h0413;
		end
		32'h00006716: begin
				q			<=			16'h0005;
		end
		32'h00006718: begin
				q			<=			16'h9597;
		end
		32'h0000671A: begin
				q			<=			16'h0000;
		end
		32'h0000671C: begin
				q			<=			16'h8593;
		end
		32'h0000671E: begin
				q			<=			16'h6985;
		end
		32'h00006720: begin
				q			<=			16'h10E3;
		end
		32'h00006722: begin
				q			<=			16'h2405;
		end
		32'h00006724: begin
				q			<=			16'h0793;
		end
		32'h00006726: begin
				q			<=			16'h0900;
		end
		32'h00006728: begin
				q			<=			16'h0593;
		end
		32'h0000672A: begin
				q			<=			16'h06C1;
		end
		32'h0000672C: begin
				q			<=			16'h0513;
		end
		32'h0000672E: begin
				q			<=			16'h0501;
		end
		32'h00006730: begin
				q			<=			16'h2A23;
		end
		32'h00006732: begin
				q			<=			16'h14F1;
		end
		32'h00006734: begin
				q			<=			16'hE0EF;
		end
		32'h00006736: begin
				q			<=			16'hAD9F;
		end
		32'h00006738: begin
				q			<=			16'h5783;
		end
		32'h0000673A: begin
				q			<=			16'h07E1;
		end
		32'h0000673C: begin
				q			<=			16'h0A93;
		end
		32'h0000673E: begin
				q			<=			16'h0000;
		end
		32'h00006740: begin
				q			<=			16'h9713;
		end
		32'h00006742: begin
				q			<=			16'h0107;
		end
		32'h00006744: begin
				q			<=			16'h5713;
		end
		32'h00006746: begin
				q			<=			16'h4107;
		end
		32'h00006748: begin
				q			<=			16'h5E63;
		end
		32'h0000674A: begin
				q			<=			16'h0007;
		end
		32'h0000674C: begin
				q			<=			16'h8737;
		end
		32'h0000674E: begin
				q			<=			16'h0000;
		end
		32'h00006750: begin
				q			<=			16'h0713;
		end
		32'h00006752: begin
				q			<=			16'hFFF7;
		end
		32'h00006754: begin
				q			<=			16'hF7B3;
		end
		32'h00006756: begin
				q			<=			16'h00E7;
		end
		32'h00006758: begin
				q			<=			16'h0AB7;
		end
		32'h0000675A: begin
				q			<=			16'h0001;
		end
		32'h0000675C: begin
				q			<=			16'h1F23;
		end
		32'h0000675E: begin
				q			<=			16'h06F1;
		end
		32'h00006760: begin
				q			<=			16'h8A93;
		end
		32'h00006762: begin
				q			<=			16'hFFFA;
		end
		32'h00006764: begin
				q			<=			16'h0593;
		end
		32'h00006766: begin
				q			<=			16'h0881;
		end
		32'h00006768: begin
				q			<=			16'h9517;
		end
		32'h0000676A: begin
				q			<=			16'h0000;
		end
		32'h0000676C: begin
				q			<=			16'h0513;
		end
		32'h0000676E: begin
				q			<=			16'hB585;
		end
		32'h00006770: begin
				q			<=			16'hE0EF;
		end
		32'h00006772: begin
				q			<=			16'hA9DF;
		end
		32'h00006774: begin
				q			<=			16'h5703;
		end
		32'h00006776: begin
				q			<=			16'h07E1;
		end
		32'h00006778: begin
				q			<=			16'h14E3;
		end
		32'h0000677A: begin
				q			<=			16'h1C07;
		end
		32'h0000677C: begin
				q			<=			16'h0713;
		end
		32'h0000677E: begin
				q			<=			16'h06C1;
		end
		32'h00006780: begin
				q			<=			16'h0793;
		end
		32'h00006782: begin
				q			<=			16'h0000;
		end
		32'h00006784: begin
				q			<=			16'h0693;
		end
		32'h00006786: begin
				q			<=			16'h0090;
		end
		32'h00006788: begin
				q			<=			16'h5603;
		end
		32'h0000678A: begin
				q			<=			16'h0007;
		end
		32'h0000678C: begin
				q			<=			16'h1A63;
		end
		32'h0000678E: begin
				q			<=			16'h1006;
		end
		32'h00006790: begin
				q			<=			16'h8793;
		end
		32'h00006792: begin
				q			<=			16'h0017;
		end
		32'h00006794: begin
				q			<=			16'h0713;
		end
		32'h00006796: begin
				q			<=			16'h0027;
		end
		32'h00006798: begin
				q			<=			16'h98E3;
		end
		32'h0000679A: begin
				q			<=			16'hFED7;
		end
		32'h0000679C: begin
				q			<=			16'h0593;
		end
		32'h0000679E: begin
				q			<=			16'h0C01;
		end
		32'h000067A0: begin
				q			<=			16'h0513;
		end
		32'h000067A2: begin
				q			<=			16'h0881;
		end
		32'h000067A4: begin
				q			<=			16'hF097;
		end
		32'h000067A6: begin
				q			<=			16'hFFFF;
		end
		32'h000067A8: begin
				q			<=			16'h80E7;
		end
		32'h000067AA: begin
				q			<=			16'hDBC0;
		end
		32'h000067AC: begin
				q			<=			16'h0593;
		end
		32'h000067AE: begin
				q			<=			16'h0881;
		end
		32'h000067B0: begin
				q			<=			16'h0513;
		end
		32'h000067B2: begin
				q			<=			16'h0C01;
		end
		32'h000067B4: begin
				q			<=			16'hE0EF;
		end
		32'h000067B6: begin
				q			<=			16'hA89F;
		end
		32'h000067B8: begin
				q			<=			16'h0593;
		end
		32'h000067BA: begin
				q			<=			16'h0C01;
		end
		32'h000067BC: begin
				q			<=			16'h0513;
		end
		32'h000067BE: begin
				q			<=			16'h06C1;
		end
		32'h000067C0: begin
				q			<=			16'hF097;
		end
		32'h000067C2: begin
				q			<=			16'hFFFF;
		end
		32'h000067C4: begin
				q			<=			16'h80E7;
		end
		32'h000067C6: begin
				q			<=			16'hDA00;
		end
		32'h000067C8: begin
				q			<=			16'h0593;
		end
		32'h000067CA: begin
				q			<=			16'h06C1;
		end
		32'h000067CC: begin
				q			<=			16'h0513;
		end
		32'h000067CE: begin
				q			<=			16'h0C01;
		end
		32'h000067D0: begin
				q			<=			16'hE0EF;
		end
		32'h000067D2: begin
				q			<=			16'hA6DF;
		end
		32'h000067D4: begin
				q			<=			16'h0613;
		end
		32'h000067D6: begin
				q			<=			16'h1501;
		end
		32'h000067D8: begin
				q			<=			16'h0593;
		end
		32'h000067DA: begin
				q			<=			16'h06C1;
		end
		32'h000067DC: begin
				q			<=			16'h0513;
		end
		32'h000067DE: begin
				q			<=			16'h0881;
		end
		32'h000067E0: begin
				q			<=			16'hF097;
		end
		32'h000067E2: begin
				q			<=			16'hFFFF;
		end
		32'h000067E4: begin
				q			<=			16'h80E7;
		end
		32'h000067E6: begin
				q			<=			16'h6E80;
		end
		32'h000067E8: begin
				q			<=			16'h5B03;
		end
		32'h000067EA: begin
				q			<=			16'h19C1;
		end
		32'h000067EC: begin
				q			<=			16'h9C17;
		end
		32'h000067EE: begin
				q			<=			16'h0000;
		end
		32'h000067F0: begin
				q			<=			16'h0C13;
		end
		32'h000067F2: begin
				q			<=			16'hAC0C;
		end
		32'h000067F4: begin
				q			<=			16'h1A63;
		end
		32'h000067F6: begin
				q			<=			16'h000B;
		end
		32'h000067F8: begin
				q			<=			16'h0593;
		end
		32'h000067FA: begin
				q			<=			16'h000C;
		end
		32'h000067FC: begin
				q			<=			16'h0513;
		end
		32'h000067FE: begin
				q			<=			16'h06C1;
		end
		32'h00006800: begin
				q			<=			16'hE0EF;
		end
		32'h00006802: begin
				q			<=			16'hE31F;
		end
		32'h00006804: begin
				q			<=			16'h1263;
		end
		32'h00006806: begin
				q			<=			16'h7005;
		end
		32'h00006808: begin
				q			<=			16'h0793;
		end
		32'h0000680A: begin
				q			<=			16'h02D0;
		end
		32'h0000680C: begin
				q			<=			16'h9463;
		end
		32'h0000680E: begin
				q			<=			16'h000A;
		end
		32'h00006810: begin
				q			<=			16'h0793;
		end
		32'h00006812: begin
				q			<=			16'h0200;
		end
		32'h00006814: begin
				q			<=			16'h0A23;
		end
		32'h00006816: begin
				q			<=			16'h10F1;
		end
		32'h00006818: begin
				q			<=			16'h0793;
		end
		32'h0000681A: begin
				q			<=			16'h0030;
		end
		32'h0000681C: begin
				q			<=			16'h8C13;
		end
		32'h0000681E: begin
				q			<=			16'h0004;
		end
		32'h00006820: begin
				q			<=			16'h1863;
		end
		32'h00006822: begin
				q			<=			16'h00FA;
		end
		32'h00006824: begin
				q			<=			16'h8C33;
		end
		32'h00006826: begin
				q			<=			16'h0084;
		end
		32'h00006828: begin
				q			<=			16'h0793;
		end
		32'h0000682A: begin
				q			<=			16'h02A0;
		end
		32'h0000682C: begin
				q			<=			16'hCAE3;
		end
		32'h0000682E: begin
				q			<=			16'h2987;
		end
		32'h00006830: begin
				q			<=			16'h0793;
		end
		32'h00006832: begin
				q			<=			16'h00A0;
		end
		32'h00006834: begin
				q			<=			16'h1863;
		end
		32'h00006836: begin
				q			<=			16'h72FB;
		end
		32'h00006838: begin
				q			<=			16'h0793;
		end
		32'h0000683A: begin
				q			<=			16'h0310;
		end
		32'h0000683C: begin
				q			<=			16'h0AA3;
		end
		32'h0000683E: begin
				q			<=			16'h10F1;
		end
		32'h00006840: begin
				q			<=			16'h0793;
		end
		32'h00006842: begin
				q			<=			16'h02E0;
		end
		32'h00006844: begin
				q			<=			16'h0B23;
		end
		32'h00006846: begin
				q			<=			16'h10F1;
		end
		32'h00006848: begin
				q			<=			16'h0B13;
		end
		32'h0000684A: begin
				q			<=			16'h1171;
		end
		32'h0000684C: begin
				q			<=			16'h5A63;
		end
		32'h0000684E: begin
				q			<=			16'h0180;
		end
		32'h00006850: begin
				q			<=			16'h0793;
		end
		32'h00006852: begin
				q			<=			16'h0300;
		end
		32'h00006854: begin
				q			<=			16'h0BA3;
		end
		32'h00006856: begin
				q			<=			16'h10F1;
		end
		32'h00006858: begin
				q			<=			16'h0C13;
		end
		32'h0000685A: begin
				q			<=			16'hFFFC;
		end
		32'h0000685C: begin
				q			<=			16'h0B13;
		end
		32'h0000685E: begin
				q			<=			16'h1181;
		end
		32'h00006860: begin
				q			<=			16'h0413;
		end
		32'h00006862: begin
				q			<=			16'h0014;
		end
		32'h00006864: begin
				q			<=			16'h5A63;
		end
		32'h00006866: begin
				q			<=			16'h700C;
		end
		32'h00006868: begin
				q			<=			16'h0613;
		end
		32'h0000686A: begin
				q			<=			16'h0004;
		end
		32'h0000686C: begin
				q			<=			16'h9597;
		end
		32'h0000686E: begin
				q			<=			16'h0000;
		end
		32'h00006870: begin
				q			<=			16'h8593;
		end
		32'h00006872: begin
				q			<=			16'h5685;
		end
		32'h00006874: begin
				q			<=			16'h0513;
		end
		32'h00006876: begin
				q			<=			16'h000B;
		end
		32'h00006878: begin
				q			<=			16'h20EF;
		end
		32'h0000687A: begin
				q			<=			16'h2440;
		end
		32'h0000687C: begin
				q			<=			16'h006F;
		end
		32'h0000687E: begin
				q			<=			16'h0F50;
		end
		32'h00006880: begin
				q			<=			16'h2023;
		end
		32'h00006882: begin
				q			<=			16'h0004;
		end
		32'h00006884: begin
				q			<=			16'hF06F;
		end
		32'h00006886: begin
				q			<=			16'hE5DF;
		end
		32'h00006888: begin
				q			<=			16'h8493;
		end
		32'h0000688A: begin
				q			<=			16'h0009;
		end
		32'h0000688C: begin
				q			<=			16'hF06F;
		end
		32'h0000688E: begin
				q			<=			16'hE69F;
		end
		32'h00006890: begin
				q			<=			16'h1783;
		end
		32'h00006892: begin
				q			<=			16'h07C1;
		end
		32'h00006894: begin
				q			<=			16'h9597;
		end
		32'h00006896: begin
				q			<=			16'h0000;
		end
		32'h00006898: begin
				q			<=			16'h8593;
		end
		32'h0000689A: begin
				q			<=			16'h53C5;
		end
		32'h0000689C: begin
				q			<=			16'hD2E3;
		end
		32'h0000689E: begin
				q			<=			16'h0C07;
		end
		32'h000068A0: begin
				q			<=			16'h0593;
		end
		32'h000068A2: begin
				q			<=			16'h06C1;
		end
		32'h000068A4: begin
				q			<=			16'h9517;
		end
		32'h000068A6: begin
				q			<=			16'h0000;
		end
		32'h000068A8: begin
				q			<=			16'h0513;
		end
		32'h000068AA: begin
				q			<=			16'hA1C5;
		end
		32'h000068AC: begin
				q			<=			16'hE0EF;
		end
		32'h000068AE: begin
				q			<=			16'hD85F;
		end
		32'h000068B0: begin
				q			<=			16'h06E3;
		end
		32'h000068B2: begin
				q			<=			16'hEE05;
		end
		32'h000068B4: begin
				q			<=			16'h5863;
		end
		32'h000068B6: begin
				q			<=			16'h4A05;
		end
		32'h000068B8: begin
				q			<=			16'h0593;
		end
		32'h000068BA: begin
				q			<=			16'h0A41;
		end
		32'h000068BC: begin
				q			<=			16'h0513;
		end
		32'h000068BE: begin
				q			<=			16'h06C1;
		end
		32'h000068C0: begin
				q			<=			16'hE0EF;
		end
		32'h000068C2: begin
				q			<=			16'h94DF;
		end
		32'h000068C4: begin
				q			<=			16'h47B7;
		end
		32'h000068C6: begin
				q			<=			16'h0000;
		end
		32'h000068C8: begin
				q			<=			16'h8793;
		end
		32'h000068CA: begin
				q			<=			16'h08E7;
		end
		32'h000068CC: begin
				q			<=			16'h1B23;
		end
		32'h000068CE: begin
				q			<=			16'h0AF1;
		end
		32'h000068D0: begin
				q			<=			16'h87B7;
		end
		32'h000068D2: begin
				q			<=			16'h0000;
		end
		32'h000068D4: begin
				q			<=			16'h8793;
		end
		32'h000068D6: begin
				q			<=			16'hFFF7;
		end
		32'h000068D8: begin
				q			<=			16'h2A23;
		end
		32'h000068DA: begin
				q			<=			16'h00F1;
		end
		32'h000068DC: begin
				q			<=			16'hC7B7;
		end
		32'h000068DE: begin
				q			<=			16'hFFFF;
		end
		32'h000068E0: begin
				q			<=			16'h8793;
		end
		32'h000068E2: begin
				q			<=			16'h0027;
		end
		32'h000068E4: begin
				q			<=			16'h0C13;
		end
		32'h000068E6: begin
				q			<=			16'h0000;
		end
		32'h000068E8: begin
				q			<=			16'h0C93;
		end
		32'h000068EA: begin
				q			<=			16'h0100;
		end
		32'h000068EC: begin
				q			<=			16'h2C23;
		end
		32'h000068EE: begin
				q			<=			16'h00F1;
		end
		32'h000068F0: begin
				q			<=			16'h9797;
		end
		32'h000068F2: begin
				q			<=			16'h0000;
		end
		32'h000068F4: begin
				q			<=			16'h8793;
		end
		32'h000068F6: begin
				q			<=			16'hA847;
		end
		32'h000068F8: begin
				q			<=			16'h8533;
		end
		32'h000068FA: begin
				q			<=			16'h0187;
		end
		32'h000068FC: begin
				q			<=			16'h0693;
		end
		32'h000068FE: begin
				q			<=			16'h1501;
		end
		32'h00006900: begin
				q			<=			16'h0613;
		end
		32'h00006902: begin
				q			<=			16'h0881;
		end
		32'h00006904: begin
				q			<=			16'h0593;
		end
		32'h00006906: begin
				q			<=			16'h0A41;
		end
		32'h00006908: begin
				q			<=			16'h0097;
		end
		32'h0000690A: begin
				q			<=			16'h0000;
		end
		32'h0000690C: begin
				q			<=			16'h80E7;
		end
		32'h0000690E: begin
				q			<=			16'h98C0;
		end
		32'h00006910: begin
				q			<=			16'h0593;
		end
		32'h00006912: begin
				q			<=			16'h03C1;
		end
		32'h00006914: begin
				q			<=			16'h0513;
		end
		32'h00006916: begin
				q			<=			16'h0881;
		end
		32'h00006918: begin
				q			<=			16'hE0EF;
		end
		32'h0000691A: begin
				q			<=			16'h8F5F;
		end
		32'h0000691C: begin
				q			<=			16'h2783;
		end
		32'h0000691E: begin
				q			<=			16'h0141;
		end
		32'h00006920: begin
				q			<=			16'h5B03;
		end
		32'h00006922: begin
				q			<=			16'h04E1;
		end
		32'h00006924: begin
				q			<=			16'h7733;
		end
		32'h00006926: begin
				q			<=			16'h00FB;
		end
		32'h00006928: begin
				q			<=			16'h2783;
		end
		32'h0000692A: begin
				q			<=			16'h0181;
		end
		32'h0000692C: begin
				q			<=			16'h0733;
		end
		32'h0000692E: begin
				q			<=			16'h00F7;
		end
		32'h00006930: begin
				q			<=			16'h4263;
		end
		32'h00006932: begin
				q			<=			16'h06E0;
		end
		32'h00006934: begin
				q			<=			16'h0513;
		end
		32'h00006936: begin
				q			<=			16'h0C01;
		end
		32'h00006938: begin
				q			<=			16'hF097;
		end
		32'h0000693A: begin
				q			<=			16'hFFFF;
		end
		32'h0000693C: begin
				q			<=			16'h80E7;
		end
		32'h0000693E: begin
				q			<=			16'h8C00;
		end
		32'h00006940: begin
				q			<=			16'h1B13;
		end
		32'h00006942: begin
				q			<=			16'h010B;
		end
		32'h00006944: begin
				q			<=			16'h5B13;
		end
		32'h00006946: begin
				q			<=			16'h410B;
		end
		32'h00006948: begin
				q			<=			16'h5A63;
		end
		32'h0000694A: begin
				q			<=			16'h120B;
		end
		32'h0000694C: begin
				q			<=			16'h0793;
		end
		32'h0000694E: begin
				q			<=			16'h0000;
		end
		32'h00006950: begin
				q			<=			16'h0713;
		end
		32'h00006952: begin
				q			<=			16'h03C1;
		end
		32'h00006954: begin
				q			<=			16'h0733;
		end
		32'h00006956: begin
				q			<=			16'h00F7;
		end
		32'h00006958: begin
				q			<=			16'h5683;
		end
		32'h0000695A: begin
				q			<=			16'h0007;
		end
		32'h0000695C: begin
				q			<=			16'h0713;
		end
		32'h0000695E: begin
				q			<=			16'h0C01;
		end
		32'h00006960: begin
				q			<=			16'h0733;
		end
		32'h00006962: begin
				q			<=			16'h00F7;
		end
		32'h00006964: begin
				q			<=			16'h5703;
		end
		32'h00006966: begin
				q			<=			16'h0007;
		end
		32'h00006968: begin
				q			<=			16'h8663;
		end
		32'h0000696A: begin
				q			<=			16'h3EE6;
		end
		32'h0000696C: begin
				q			<=			16'h9517;
		end
		32'h0000696E: begin
				q			<=			16'h0000;
		end
		32'h00006970: begin
				q			<=			16'h0513;
		end
		32'h00006972: begin
				q			<=			16'h9545;
		end
		32'h00006974: begin
				q			<=			16'hF097;
		end
		32'h00006976: begin
				q			<=			16'hFFFF;
		end
		32'h00006978: begin
				q			<=			16'h80E7;
		end
		32'h0000697A: begin
				q			<=			16'hB7C0;
		end
		32'h0000697C: begin
				q			<=			16'h0863;
		end
		32'h0000697E: begin
				q			<=			16'h0805;
		end
		32'h00006980: begin
				q			<=			16'h0593;
		end
		32'h00006982: begin
				q			<=			16'h0C01;
		end
		32'h00006984: begin
				q			<=			16'h9517;
		end
		32'h00006986: begin
				q			<=			16'h0000;
		end
		32'h00006988: begin
				q			<=			16'h0513;
		end
		32'h0000698A: begin
				q			<=			16'h93C5;
		end
		32'h0000698C: begin
				q			<=			16'hE0EF;
		end
		32'h0000698E: begin
				q			<=			16'h881F;
		end
		32'h00006990: begin
				q			<=			16'h006F;
		end
		32'h00006992: begin
				q			<=			16'h0EC0;
		end
		32'h00006994: begin
				q			<=			16'h0793;
		end
		32'h00006996: begin
				q			<=			16'h0900;
		end
		32'h00006998: begin
				q			<=			16'h8D33;
		end
		32'h0000699A: begin
				q			<=			16'h40E7;
		end
		32'h0000699C: begin
				q			<=			16'h0593;
		end
		32'h0000699E: begin
				q			<=			16'h0C01;
		end
		32'h000069A0: begin
				q			<=			16'h0513;
		end
		32'h000069A2: begin
				q			<=			16'h03C1;
		end
		32'h000069A4: begin
				q			<=			16'hE0EF;
		end
		32'h000069A6: begin
				q			<=			16'h869F;
		end
		32'h000069A8: begin
				q			<=			16'h5A63;
		end
		32'h000069AA: begin
				q			<=			16'h0DA0;
		end
		32'h000069AC: begin
				q			<=			16'h0693;
		end
		32'h000069AE: begin
				q			<=			16'h0C01;
		end
		32'h000069B0: begin
				q			<=			16'h0793;
		end
		32'h000069B2: begin
				q			<=			16'h000D;
		end
		32'h000069B4: begin
				q			<=			16'h0613;
		end
		32'h000069B6: begin
				q			<=			16'h00F0;
		end
		32'h000069B8: begin
				q			<=			16'h4263;
		end
		32'h000069BA: begin
				q			<=			16'h04F6;
		end
		32'h000069BC: begin
				q			<=			16'h5793;
		end
		32'h000069BE: begin
				q			<=			16'h004D;
		end
		32'h000069C0: begin
				q			<=			16'h0613;
		end
		32'h000069C2: begin
				q			<=			16'hFF00;
		end
		32'h000069C4: begin
				q			<=			16'h9693;
		end
		32'h000069C6: begin
				q			<=			16'h0017;
		end
		32'h000069C8: begin
				q			<=			16'h87B3;
		end
		32'h000069CA: begin
				q			<=			16'h02C7;
		end
		32'h000069CC: begin
				q			<=			16'h0713;
		end
		32'h000069CE: begin
				q			<=			16'h0C01;
		end
		32'h000069D0: begin
				q			<=			16'h06B3;
		end
		32'h000069D2: begin
				q			<=			16'h00D7;
		end
		32'h000069D4: begin
				q			<=			16'h9717;
		end
		32'h000069D6: begin
				q			<=			16'h0000;
		end
		32'h000069D8: begin
				q			<=			16'h0713;
		end
		32'h000069DA: begin
				q			<=			16'h8D87;
		end
		32'h000069DC: begin
				q			<=			16'h87B3;
		end
		32'h000069DE: begin
				q			<=			16'h01A7;
		end
		32'h000069E0: begin
				q			<=			16'h9793;
		end
		32'h000069E2: begin
				q			<=			16'h0017;
		end
		32'h000069E4: begin
				q			<=			16'h07B3;
		end
		32'h000069E6: begin
				q			<=			16'h00F7;
		end
		32'h000069E8: begin
				q			<=			16'hD783;
		end
		32'h000069EA: begin
				q			<=			16'h12C7;
		end
		32'h000069EC: begin
				q			<=			16'hD703;
		end
		32'h000069EE: begin
				q			<=			16'h0006;
		end
		32'h000069F0: begin
				q			<=			16'hF7B3;
		end
		32'h000069F2: begin
				q			<=			16'h00E7;
		end
		32'h000069F4: begin
				q			<=			16'h9023;
		end
		32'h000069F6: begin
				q			<=			16'h00F6;
		end
		32'h000069F8: begin
				q			<=			16'hF06F;
		end
		32'h000069FA: begin
				q			<=			16'hF49F;
		end
		32'h000069FC: begin
				q			<=			16'h9023;
		end
		32'h000069FE: begin
				q			<=			16'h0006;
		end
		32'h00006A00: begin
				q			<=			16'h8793;
		end
		32'h00006A02: begin
				q			<=			16'hFF07;
		end
		32'h00006A04: begin
				q			<=			16'h8693;
		end
		32'h00006A06: begin
				q			<=			16'h0026;
		end
		32'h00006A08: begin
				q			<=			16'hF06F;
		end
		32'h00006A0A: begin
				q			<=			16'hFB1F;
		end
		32'h00006A0C: begin
				q			<=			16'h0513;
		end
		32'h00006A0E: begin
				q			<=			16'h0C01;
		end
		32'h00006A10: begin
				q			<=			16'hF097;
		end
		32'h00006A12: begin
				q			<=			16'hFFFF;
		end
		32'h00006A14: begin
				q			<=			16'h80E7;
		end
		32'h00006A16: begin
				q			<=			16'hAE00;
		end
		32'h00006A18: begin
				q			<=			16'h0863;
		end
		32'h00006A1A: begin
				q			<=			16'h0005;
		end
		32'h00006A1C: begin
				q			<=			16'h0593;
		end
		32'h00006A1E: begin
				q			<=			16'h0C01;
		end
		32'h00006A20: begin
				q			<=			16'h8513;
		end
		32'h00006A22: begin
				q			<=			16'h0005;
		end
		32'h00006A24: begin
				q			<=			16'hF06F;
		end
		32'h00006A26: begin
				q			<=			16'hF69F;
		end
		32'h00006A28: begin
				q			<=			16'h9517;
		end
		32'h00006A2A: begin
				q			<=			16'h0000;
		end
		32'h00006A2C: begin
				q			<=			16'h0513;
		end
		32'h00006A2E: begin
				q			<=			16'h8985;
		end
		32'h00006A30: begin
				q			<=			16'hF097;
		end
		32'h00006A32: begin
				q			<=			16'hFFFF;
		end
		32'h00006A34: begin
				q			<=			16'h80E7;
		end
		32'h00006A36: begin
				q			<=			16'hD180;
		end
		32'h00006A38: begin
				q			<=			16'h0D13;
		end
		32'h00006A3A: begin
				q			<=			16'h0005;
		end
		32'h00006A3C: begin
				q			<=			16'h0513;
		end
		32'h00006A3E: begin
				q			<=			16'h0C01;
		end
		32'h00006A40: begin
				q			<=			16'hF097;
		end
		32'h00006A42: begin
				q			<=			16'hFFFF;
		end
		32'h00006A44: begin
				q			<=			16'h80E7;
		end
		32'h00006A46: begin
				q			<=			16'hD080;
		end
		32'h00006A48: begin
				q			<=			16'h0B13;
		end
		32'h00006A4A: begin
				q			<=			16'h0005;
		end
		32'h00006A4C: begin
				q			<=			16'h0263;
		end
		32'h00006A4E: begin
				q			<=			16'h160D;
		end
		32'h00006A50: begin
				q			<=			16'h0663;
		end
		32'h00006A52: begin
				q			<=			16'h1205;
		end
		32'h00006A54: begin
				q			<=			16'h9517;
		end
		32'h00006A56: begin
				q			<=			16'h0000;
		end
		32'h00006A58: begin
				q			<=			16'h0513;
		end
		32'h00006A5A: begin
				q			<=			16'h86C5;
		end
		32'h00006A5C: begin
				q			<=			16'hE0EF;
		end
		32'h00006A5E: begin
				q			<=			16'hAC9F;
		end
		32'h00006A60: begin
				q			<=			16'h0B13;
		end
		32'h00006A62: begin
				q			<=			16'h0005;
		end
		32'h00006A64: begin
				q			<=			16'h0513;
		end
		32'h00006A66: begin
				q			<=			16'h0C01;
		end
		32'h00006A68: begin
				q			<=			16'hE0EF;
		end
		32'h00006A6A: begin
				q			<=			16'hABDF;
		end
		32'h00006A6C: begin
				q			<=			16'h1863;
		end
		32'h00006A6E: begin
				q			<=			16'h10AB;
		end
		32'h00006A70: begin
				q			<=			16'h0513;
		end
		32'h00006A72: begin
				q			<=			16'h0C01;
		end
		32'h00006A74: begin
				q			<=			16'hF097;
		end
		32'h00006A76: begin
				q			<=			16'hFFFF;
		end
		32'h00006A78: begin
				q			<=			16'h80E7;
		end
		32'h00006A7A: begin
				q			<=			16'hF740;
		end
		32'h00006A7C: begin
				q			<=			16'h0793;
		end
		32'h00006A7E: begin
				q			<=			16'h0000;
		end
		32'h00006A80: begin
				q			<=			16'h0713;
		end
		32'h00006A82: begin
				q			<=			16'h0881;
		end
		32'h00006A84: begin
				q			<=			16'h0733;
		end
		32'h00006A86: begin
				q			<=			16'h00F7;
		end
		32'h00006A88: begin
				q			<=			16'h5683;
		end
		32'h00006A8A: begin
				q			<=			16'h0007;
		end
		32'h00006A8C: begin
				q			<=			16'h0713;
		end
		32'h00006A8E: begin
				q			<=			16'h0C01;
		end
		32'h00006A90: begin
				q			<=			16'h0733;
		end
		32'h00006A92: begin
				q			<=			16'h00F7;
		end
		32'h00006A94: begin
				q			<=			16'h5703;
		end
		32'h00006A96: begin
				q			<=			16'h0007;
		end
		32'h00006A98: begin
				q			<=			16'h9063;
		end
		32'h00006A9A: begin
				q			<=			16'h02E6;
		end
		32'h00006A9C: begin
				q			<=			16'h8793;
		end
		32'h00006A9E: begin
				q			<=			16'h0027;
		end
		32'h00006AA0: begin
				q			<=			16'h0713;
		end
		32'h00006AA2: begin
				q			<=			16'h0120;
		end
		32'h00006AA4: begin
				q			<=			16'h9EE3;
		end
		32'h00006AA6: begin
				q			<=			16'hFCE7;
		end
		32'h00006AA8: begin
				q			<=			16'h0593;
		end
		32'h00006AAA: begin
				q			<=			16'h0A41;
		end
		32'h00006AAC: begin
				q			<=			16'h0513;
		end
		32'h00006AAE: begin
				q			<=			16'h0881;
		end
		32'h00006AB0: begin
				q			<=			16'hE0EF;
		end
		32'h00006AB2: begin
				q			<=			16'hF5CF;
		end
		32'h00006AB4: begin
				q			<=			16'h0433;
		end
		32'h00006AB6: begin
				q			<=			16'h0194;
		end
		32'h00006AB8: begin
				q			<=			16'h0C13;
		end
		32'h00006ABA: begin
				q			<=			16'h014C;
		end
		32'h00006ABC: begin
				q			<=			16'h0793;
		end
		32'h00006ABE: begin
				q			<=			16'h0640;
		end
		32'h00006AC0: begin
				q			<=			16'hDC93;
		end
		32'h00006AC2: begin
				q			<=			16'h001C;
		end
		32'h00006AC4: begin
				q			<=			16'h16E3;
		end
		32'h00006AC6: begin
				q			<=			16'hE2FC;
		end
		32'h00006AC8: begin
				q			<=			16'h5783;
		end
		32'h00006ACA: begin
				q			<=			16'h0B61;
		end
		32'h00006ACC: begin
				q			<=			16'h5703;
		end
		32'h00006ACE: begin
				q			<=			16'h07E1;
		end
		32'h00006AD0: begin
				q			<=			16'h0593;
		end
		32'h00006AD2: begin
				q			<=			16'h06C1;
		end
		32'h00006AD4: begin
				q			<=			16'h0513;
		end
		32'h00006AD6: begin
				q			<=			16'h0A41;
		end
		32'h00006AD8: begin
				q			<=			16'h87B3;
		end
		32'h00006ADA: begin
				q			<=			16'h00E7;
		end
		32'h00006ADC: begin
				q			<=			16'hC737;
		end
		32'h00006ADE: begin
				q			<=			16'hFFFF;
		end
		32'h00006AE0: begin
				q			<=			16'h0713;
		end
		32'h00006AE2: begin
				q			<=			16'hF727;
		end
		32'h00006AE4: begin
				q			<=			16'h87B3;
		end
		32'h00006AE6: begin
				q			<=			16'h00E7;
		end
		32'h00006AE8: begin
				q			<=			16'h1B23;
		end
		32'h00006AEA: begin
				q			<=			16'h0AF1;
		end
		32'h00006AEC: begin
				q			<=			16'hE0EF;
		end
		32'h00006AEE: begin
				q			<=			16'hF20F;
		end
		32'h00006AF0: begin
				q			<=			16'h0593;
		end
		32'h00006AF2: begin
				q			<=			16'h0881;
		end
		32'h00006AF4: begin
				q			<=			16'h8517;
		end
		32'h00006AF6: begin
				q			<=			16'h0000;
		end
		32'h00006AF8: begin
				q			<=			16'h0513;
		end
		32'h00006AFA: begin
				q			<=			16'h7CC5;
		end
		32'h00006AFC: begin
				q			<=			16'hE0EF;
		end
		32'h00006AFE: begin
				q			<=			16'hF10F;
		end
		32'h00006B00: begin
				q			<=			16'h0B13;
		end
		32'h00006B02: begin
				q			<=			16'h0000;
		end
		32'h00006B04: begin
				q			<=			16'h1CB7;
		end
		32'h00006B06: begin
				q			<=			16'h0000;
		end
		32'h00006B08: begin
				q			<=			16'h0D93;
		end
		32'h00006B0A: begin
				q			<=			16'h1040;
		end
		32'h00006B0C: begin
				q			<=			16'h8797;
		end
		32'h00006B0E: begin
				q			<=			16'h0000;
		end
		32'h00006B10: begin
				q			<=			16'h8793;
		end
		32'h00006B12: begin
				q			<=			16'h7C87;
		end
		32'h00006B14: begin
				q			<=			16'h0593;
		end
		32'h00006B16: begin
				q			<=			16'h0A41;
		end
		32'h00006B18: begin
				q			<=			16'h9517;
		end
		32'h00006B1A: begin
				q			<=			16'h0000;
		end
		32'h00006B1C: begin
				q			<=			16'h0513;
		end
		32'h00006B1E: begin
				q			<=			16'h8AC5;
		end
		32'h00006B20: begin
				q			<=			16'h0C33;
		end
		32'h00006B22: begin
				q			<=			16'h00FB;
		end
		32'h00006B24: begin
				q			<=			16'hE0EF;
		end
		32'h00006B26: begin
				q			<=			16'hB0DF;
		end
		32'h00006B28: begin
				q			<=			16'h4AE3;
		end
		32'h00006B2A: begin
				q			<=			16'hC6A0;
		end
		32'h00006B2C: begin
				q			<=			16'h0593;
		end
		32'h00006B2E: begin
				q			<=			16'h0A41;
		end
		32'h00006B30: begin
				q			<=			16'h0513;
		end
		32'h00006B32: begin
				q			<=			16'h000C;
		end
		32'h00006B34: begin
				q			<=			16'hE0EF;
		end
		32'h00006B36: begin
				q			<=			16'hAFDF;
		end
		32'h00006B38: begin
				q			<=			16'h4A63;
		end
		32'h00006B3A: begin
				q			<=			16'h02A0;
		end
		32'h00006B3C: begin
				q			<=			16'h0613;
		end
		32'h00006B3E: begin
				q			<=			16'h0A41;
		end
		32'h00006B40: begin
				q			<=			16'h0593;
		end
		32'h00006B42: begin
				q			<=			16'h0006;
		end
		32'h00006B44: begin
				q			<=			16'h0693;
		end
		32'h00006B46: begin
				q			<=			16'h1501;
		end
		32'h00006B48: begin
				q			<=			16'h0513;
		end
		32'h00006B4A: begin
				q			<=			16'h000C;
		end
		32'h00006B4C: begin
				q			<=			16'hF097;
		end
		32'h00006B4E: begin
				q			<=			16'hFFFF;
		end
		32'h00006B50: begin
				q			<=			16'h80E7;
		end
		32'h00006B52: begin
				q			<=			16'h7480;
		end
		32'h00006B54: begin
				q			<=			16'h0613;
		end
		32'h00006B56: begin
				q			<=			16'h0881;
		end
		32'h00006B58: begin
				q			<=			16'h0693;
		end
		32'h00006B5A: begin
				q			<=			16'h1501;
		end
		32'h00006B5C: begin
				q			<=			16'h0593;
		end
		32'h00006B5E: begin
				q			<=			16'h0006;
		end
		32'h00006B60: begin
				q			<=			16'h0513;
		end
		32'h00006B62: begin
				q			<=			16'h000C;
		end
		32'h00006B64: begin
				q			<=			16'hF0EF;
		end
		32'h00006B66: begin
				q			<=			16'hC54F;
		end
		32'h00006B68: begin
				q			<=			16'h0433;
		end
		32'h00006B6A: begin
				q			<=			16'h0194;
		end
		32'h00006B6C: begin
				q			<=			16'h0B13;
		end
		32'h00006B6E: begin
				q			<=			16'h014B;
		end
		32'h00006B70: begin
				q			<=			16'hDC93;
		end
		32'h00006B72: begin
				q			<=			16'h001C;
		end
		32'h00006B74: begin
				q			<=			16'h1CE3;
		end
		32'h00006B76: begin
				q			<=			16'hF9BB;
		end
		32'h00006B78: begin
				q			<=			16'hF06F;
		end
		32'h00006B7A: begin
				q			<=			16'hC25F;
		end
		32'h00006B7C: begin
				q			<=			16'h8517;
		end
		32'h00006B7E: begin
				q			<=			16'h0000;
		end
		32'h00006B80: begin
				q			<=			16'h0513;
		end
		32'h00006B82: begin
				q			<=			16'h7445;
		end
		32'h00006B84: begin
				q			<=			16'h0593;
		end
		32'h00006B86: begin
				q			<=			16'h0C01;
		end
		32'h00006B88: begin
				q			<=			16'hE0EF;
		end
		32'h00006B8A: begin
				q			<=			16'hE84F;
		end
		32'h00006B8C: begin
				q			<=			16'h0513;
		end
		32'h00006B8E: begin
				q			<=			16'h0C01;
		end
		32'h00006B90: begin
				q			<=			16'hF097;
		end
		32'h00006B92: begin
				q			<=			16'hFFFF;
		end
		32'h00006B94: begin
				q			<=			16'h80E7;
		end
		32'h00006B96: begin
				q			<=			16'h9600;
		end
		32'h00006B98: begin
				q			<=			16'h12E3;
		end
		32'h00006B9A: begin
				q			<=			16'hEE05;
		end
		32'h00006B9C: begin
				q			<=			16'h5783;
		end
		32'h00006B9E: begin
				q			<=			16'h0D21;
		end
		32'h00006BA0: begin
				q			<=			16'h8737;
		end
		32'h00006BA2: begin
				q			<=			16'hFFFF;
		end
		32'h00006BA4: begin
				q			<=			16'hC7B3;
		end
		32'h00006BA6: begin
				q			<=			16'h00E7;
		end
		32'h00006BA8: begin
				q			<=			16'h1923;
		end
		32'h00006BAA: begin
				q			<=			16'h0CF1;
		end
		32'h00006BAC: begin
				q			<=			16'hF06F;
		end
		32'h00006BAE: begin
				q			<=			16'hED1F;
		end
		32'h00006BB0: begin
				q			<=			16'h16E3;
		end
		32'h00006BB2: begin
				q			<=			16'hE605;
		end
		32'h00006BB4: begin
				q			<=			16'h0593;
		end
		32'h00006BB6: begin
				q			<=			16'h0DC1;
		end
		32'h00006BB8: begin
				q			<=			16'h8517;
		end
		32'h00006BBA: begin
				q			<=			16'h0000;
		end
		32'h00006BBC: begin
				q			<=			16'h0513;
		end
		32'h00006BBE: begin
				q			<=			16'h7085;
		end
		32'h00006BC0: begin
				q			<=			16'hF097;
		end
		32'h00006BC2: begin
				q			<=			16'hFFFF;
		end
		32'h00006BC4: begin
				q			<=			16'h80E7;
		end
		32'h00006BC6: begin
				q			<=			16'h9A00;
		end
		32'h00006BC8: begin
				q			<=			16'h0593;
		end
		32'h00006BCA: begin
				q			<=			16'h0F81;
		end
		32'h00006BCC: begin
				q			<=			16'h0513;
		end
		32'h00006BCE: begin
				q			<=			16'h0C01;
		end
		32'h00006BD0: begin
				q			<=			16'hF097;
		end
		32'h00006BD2: begin
				q			<=			16'hFFFF;
		end
		32'h00006BD4: begin
				q			<=			16'h80E7;
		end
		32'h00006BD6: begin
				q			<=			16'h9900;
		end
		32'h00006BD8: begin
				q			<=			16'h5703;
		end
		32'h00006BDA: begin
				q			<=			16'h0DC1;
		end
		32'h00006BDC: begin
				q			<=			16'h5D83;
		end
		32'h00006BDE: begin
				q			<=			16'h0FA1;
		end
		32'h00006BE0: begin
				q			<=			16'h5783;
		end
		32'h00006BE2: begin
				q			<=			16'h0DE1;
		end
		32'h00006BE4: begin
				q			<=			16'h4713;
		end
		32'h00006BE6: begin
				q			<=			16'hFFF7;
		end
		32'h00006BE8: begin
				q			<=			16'h1D13;
		end
		32'h00006BEA: begin
				q			<=			16'h0107;
		end
		32'h00006BEC: begin
				q			<=			16'h5D13;
		end
		32'h00006BEE: begin
				q			<=			16'h010D;
		end
		32'h00006BF0: begin
				q			<=			16'h1E23;
		end
		32'h00006BF2: begin
				q			<=			16'h0DA1;
		end
		32'h00006BF4: begin
				q			<=			16'h87B3;
		end
		32'h00006BF6: begin
				q			<=			16'h41B7;
		end
		32'h00006BF8: begin
				q			<=			16'h5663;
		end
		32'h00006BFA: begin
				q			<=			16'h08F0;
		end
		32'h00006BFC: begin
				q			<=			16'h0593;
		end
		32'h00006BFE: begin
				q			<=			16'h1141;
		end
		32'h00006C00: begin
				q			<=			16'h0513;
		end
		32'h00006C02: begin
				q			<=			16'h0F81;
		end
		32'h00006C04: begin
				q			<=			16'h2E23;
		end
		32'h00006C06: begin
				q			<=			16'h00F1;
		end
		32'h00006C08: begin
				q			<=			16'hE0EF;
		end
		32'h00006C0A: begin
				q			<=			16'hE34F;
		end
		32'h00006C0C: begin
				q			<=			16'h0593;
		end
		32'h00006C0E: begin
				q			<=			16'h0F81;
		end
		32'h00006C10: begin
				q			<=			16'h0513;
		end
		32'h00006C12: begin
				q			<=			16'h0DC1;
		end
		32'h00006C14: begin
				q			<=			16'hE0EF;
		end
		32'h00006C16: begin
				q			<=			16'hE28F;
		end
		32'h00006C18: begin
				q			<=			16'h0593;
		end
		32'h00006C1A: begin
				q			<=			16'h0DC1;
		end
		32'h00006C1C: begin
				q			<=			16'h0513;
		end
		32'h00006C1E: begin
				q			<=			16'h1141;
		end
		32'h00006C20: begin
				q			<=			16'hE0EF;
		end
		32'h00006C22: begin
				q			<=			16'hE1CF;
		end
		32'h00006C24: begin
				q			<=			16'h2783;
		end
		32'h00006C26: begin
				q			<=			16'h01C1;
		end
		32'h00006C28: begin
				q			<=			16'h5D83;
		end
		32'h00006C2A: begin
				q			<=			16'h0FA1;
		end
		32'h00006C2C: begin
				q			<=			16'h07B3;
		end
		32'h00006C2E: begin
				q			<=			16'h40F0;
		end
		32'h00006C30: begin
				q			<=			16'h0713;
		end
		32'h00006C32: begin
				q			<=			16'hF6F0;
		end
		32'h00006C34: begin
				q			<=			16'hCE63;
		end
		32'h00006C36: begin
				q			<=			16'h08E7;
		end
		32'h00006C38: begin
				q			<=			16'h8593;
		end
		32'h00006C3A: begin
				q			<=			16'h0007;
		end
		32'h00006C3C: begin
				q			<=			16'h0513;
		end
		32'h00006C3E: begin
				q			<=			16'h0DC1;
		end
		32'h00006C40: begin
				q			<=			16'hF097;
		end
		32'h00006C42: begin
				q			<=			16'hFFFF;
		end
		32'h00006C44: begin
				q			<=			16'h80E7;
		end
		32'h00006C46: begin
				q			<=			16'hB640;
		end
		32'h00006C48: begin
				q			<=			16'h0D13;
		end
		32'h00006C4A: begin
				q			<=			16'h0005;
		end
		32'h00006C4C: begin
				q			<=			16'h5703;
		end
		32'h00006C4E: begin
				q			<=			16'h0DC1;
		end
		32'h00006C50: begin
				q			<=			16'h5783;
		end
		32'h00006C52: begin
				q			<=			16'h0F81;
		end
		32'h00006C54: begin
				q			<=			16'h0593;
		end
		32'h00006C56: begin
				q			<=			16'h0F81;
		end
		32'h00006C58: begin
				q			<=			16'h0513;
		end
		32'h00006C5A: begin
				q			<=			16'h0DC1;
		end
		32'h00006C5C: begin
				q			<=			16'h1463;
		end
		32'h00006C5E: begin
				q			<=			16'h0EF7;
		end
		32'h00006C60: begin
				q			<=			16'hE0EF;
		end
		32'h00006C62: begin
				q			<=			16'hF84F;
		end
		32'h00006C64: begin
				q			<=			16'h0793;
		end
		32'h00006C66: begin
				q			<=			16'h1501;
		end
		32'h00006C68: begin
				q			<=			16'h0713;
		end
		32'h00006C6A: begin
				q			<=			16'h0400;
		end
		32'h00006C6C: begin
				q			<=			16'h8693;
		end
		32'h00006C6E: begin
				q			<=			16'h000D;
		end
		32'h00006C70: begin
				q			<=			16'h0613;
		end
		32'h00006C72: begin
				q			<=			16'h000B;
		end
		32'h00006C74: begin
				q			<=			16'h0593;
		end
		32'h00006C76: begin
				q			<=			16'h000D;
		end
		32'h00006C78: begin
				q			<=			16'h0513;
		end
		32'h00006C7A: begin
				q			<=			16'h0F81;
		end
		32'h00006C7C: begin
				q			<=			16'hE0EF;
		end
		32'h00006C7E: begin
				q			<=			16'hF19F;
		end
		32'h00006C80: begin
				q			<=			16'h006F;
		end
		32'h00006C82: begin
				q			<=			16'h0500;
		end
		32'h00006C84: begin
				q			<=			16'h96E3;
		end
		32'h00006C86: begin
				q			<=			16'hFA07;
		end
		32'h00006C88: begin
				q			<=			16'h0593;
		end
		32'h00006C8A: begin
				q			<=			16'h0F81;
		end
		32'h00006C8C: begin
				q			<=			16'h0513;
		end
		32'h00006C8E: begin
				q			<=			16'h0DC1;
		end
		32'h00006C90: begin
				q			<=			16'hE097;
		end
		32'h00006C92: begin
				q			<=			16'hFFFF;
		end
		32'h00006C94: begin
				q			<=			16'h80E7;
		end
		32'h00006C96: begin
				q			<=			16'h5D00;
		end
		32'h00006C98: begin
				q			<=			16'h1C63;
		end
		32'h00006C9A: begin
				q			<=			16'h0605;
		end
		32'h00006C9C: begin
				q			<=			16'h5783;
		end
		32'h00006C9E: begin
				q			<=			16'h0F81;
		end
		32'h00006CA0: begin
				q			<=			16'h8A63;
		end
		32'h00006CA2: begin
				q			<=			16'h01A7;
		end
		32'h00006CA4: begin
				q			<=			16'h0513;
		end
		32'h00006CA6: begin
				q			<=			16'h0C01;
		end
		32'h00006CA8: begin
				q			<=			16'hE097;
		end
		32'h00006CAA: begin
				q			<=			16'hFFFF;
		end
		32'h00006CAC: begin
				q			<=			16'h80E7;
		end
		32'h00006CAE: begin
				q			<=			16'h5500;
		end
		32'h00006CB0: begin
				q			<=			16'hF06F;
		end
		32'h00006CB2: begin
				q			<=			16'hDCDF;
		end
		32'h00006CB4: begin
				q			<=			16'h9663;
		end
		32'h00006CB6: begin
				q			<=			16'h020D;
		end
		32'h00006CB8: begin
				q			<=			16'h1703;
		end
		32'h00006CBA: begin
				q			<=			16'h0FE1;
		end
		32'h00006CBC: begin
				q			<=			16'h0793;
		end
		32'h00006CBE: begin
				q			<=			16'h0000;
		end
		32'h00006CC0: begin
				q			<=			16'h4263;
		end
		32'h00006CC2: begin
				q			<=			16'h0207;
		end
		32'h00006CC4: begin
				q			<=			16'h0513;
		end
		32'h00006CC6: begin
				q			<=			16'h0F81;
		end
		32'h00006CC8: begin
				q			<=			16'hE097;
		end
		32'h00006CCA: begin
				q			<=			16'hFFFF;
		end
		32'h00006CCC: begin
				q			<=			16'h80E7;
		end
		32'h00006CCE: begin
				q			<=			16'h6240;
		end
		32'h00006CD0: begin
				q			<=			16'h0593;
		end
		32'h00006CD2: begin
				q			<=			16'h0C01;
		end
		32'h00006CD4: begin
				q			<=			16'h0513;
		end
		32'h00006CD6: begin
				q			<=			16'h0F81;
		end
		32'h00006CD8: begin
				q			<=			16'hE0EF;
		end
		32'h00006CDA: begin
				q			<=			16'hD39F;
		end
		32'h00006CDC: begin
				q			<=			16'hF06F;
		end
		32'h00006CDE: begin
				q			<=			16'hDA1F;
		end
		32'h00006CE0: begin
				q			<=			16'h0793;
		end
		32'h00006CE2: begin
				q			<=			16'h0000;
		end
		32'h00006CE4: begin
				q			<=			16'h0713;
		end
		32'h00006CE6: begin
				q			<=			16'h0160;
		end
		32'h00006CE8: begin
				q			<=			16'h0693;
		end
		32'h00006CEA: begin
				q			<=			16'h0F81;
		end
		32'h00006CEC: begin
				q			<=			16'h8633;
		end
		32'h00006CEE: begin
				q			<=			16'h00F6;
		end
		32'h00006CF0: begin
				q			<=			16'h5603;
		end
		32'h00006CF2: begin
				q			<=			16'h0026;
		end
		32'h00006CF4: begin
				q			<=			16'h0863;
		end
		32'h00006CF6: begin
				q			<=			16'h0006;
		end
		32'h00006CF8: begin
				q			<=			16'h8D93;
		end
		32'h00006CFA: begin
				q			<=			16'h001D;
		end
		32'h00006CFC: begin
				q			<=			16'h1D23;
		end
		32'h00006CFE: begin
				q			<=			16'h0FB1;
		end
		32'h00006D00: begin
				q			<=			16'hF06F;
		end
		32'h00006D02: begin
				q			<=			16'hFD1F;
		end
		32'h00006D04: begin
				q			<=			16'h8793;
		end
		32'h00006D06: begin
				q			<=			16'h0027;
		end
		32'h00006D08: begin
				q			<=			16'h90E3;
		end
		32'h00006D0A: begin
				q			<=			16'hFEE7;
		end
		32'h00006D0C: begin
				q			<=			16'hF06F;
		end
		32'h00006D0E: begin
				q			<=			16'hFF1F;
		end
		32'h00006D10: begin
				q			<=			16'h0D13;
		end
		32'h00006D12: begin
				q			<=			16'h0000;
		end
		32'h00006D14: begin
				q			<=			16'h5CE3;
		end
		32'h00006D16: begin
				q			<=			16'hF2A0;
		end
		32'h00006D18: begin
				q			<=			16'h0593;
		end
		32'h00006D1A: begin
				q			<=			16'h1141;
		end
		32'h00006D1C: begin
				q			<=			16'h0513;
		end
		32'h00006D1E: begin
				q			<=			16'h0F81;
		end
		32'h00006D20: begin
				q			<=			16'hE0EF;
		end
		32'h00006D22: begin
				q			<=			16'hD1CF;
		end
		32'h00006D24: begin
				q			<=			16'h0593;
		end
		32'h00006D26: begin
				q			<=			16'h0F81;
		end
		32'h00006D28: begin
				q			<=			16'h0513;
		end
		32'h00006D2A: begin
				q			<=			16'h0DC1;
		end
		32'h00006D2C: begin
				q			<=			16'hE0EF;
		end
		32'h00006D2E: begin
				q			<=			16'hD10F;
		end
		32'h00006D30: begin
				q			<=			16'h0593;
		end
		32'h00006D32: begin
				q			<=			16'h0DC1;
		end
		32'h00006D34: begin
				q			<=			16'h0513;
		end
		32'h00006D36: begin
				q			<=			16'h1141;
		end
		32'h00006D38: begin
				q			<=			16'hE0EF;
		end
		32'h00006D3A: begin
				q			<=			16'hD04F;
		end
		32'h00006D3C: begin
				q			<=			16'h0D13;
		end
		32'h00006D3E: begin
				q			<=			16'h000B;
		end
		32'h00006D40: begin
				q			<=			16'hF06F;
		end
		32'h00006D42: begin
				q			<=			16'hF0DF;
		end
		32'h00006D44: begin
				q			<=			16'hE097;
		end
		32'h00006D46: begin
				q			<=			16'hFFFF;
		end
		32'h00006D48: begin
				q			<=			16'h80E7;
		end
		32'h00006D4A: begin
				q			<=			16'h6D80;
		end
		32'h00006D4C: begin
				q			<=			16'h0B13;
		end
		32'h00006D4E: begin
				q			<=			16'h0010;
		end
		32'h00006D50: begin
				q			<=			16'hF06F;
		end
		32'h00006D52: begin
				q			<=			16'hF15F;
		end
		32'h00006D54: begin
				q			<=			16'h8793;
		end
		32'h00006D56: begin
				q			<=			16'h0027;
		end
		32'h00006D58: begin
				q			<=			16'h0713;
		end
		32'h00006D5A: begin
				q			<=			16'h0120;
		end
		32'h00006D5C: begin
				q			<=			16'h9AE3;
		end
		32'h00006D5E: begin
				q			<=			16'hBEE7;
		end
		32'h00006D60: begin
				q			<=			16'hF06F;
		end
		32'h00006D62: begin
				q			<=			16'hD1DF;
		end
		32'h00006D64: begin
				q			<=			16'h5783;
		end
		32'h00006D66: begin
				q			<=			16'h07E1;
		end
		32'h00006D68: begin
				q			<=			16'h8B17;
		end
		32'h00006D6A: begin
				q			<=			16'h0000;
		end
		32'h00006D6C: begin
				q			<=			16'h0B13;
		end
		32'h00006D6E: begin
				q			<=			16'h65CB;
		end
		32'h00006D70: begin
				q			<=			16'h8A63;
		end
		32'h00006D72: begin
				q			<=			16'h0A07;
		end
		32'h00006D74: begin
				q			<=			16'h0593;
		end
		32'h00006D76: begin
				q			<=			16'h0C01;
		end
		32'h00006D78: begin
				q			<=			16'h0513;
		end
		32'h00006D7A: begin
				q			<=			16'h06C1;
		end
		32'h00006D7C: begin
				q			<=			16'h4B37;
		end
		32'h00006D7E: begin
				q			<=			16'h0000;
		end
		32'h00006D80: begin
				q			<=			16'hE097;
		end
		32'h00006D82: begin
				q			<=			16'hFFFF;
		end
		32'h00006D84: begin
				q			<=			16'h80E7;
		end
		32'h00006D86: begin
				q			<=			16'h7E00;
		end
		32'h00006D88: begin
				q			<=			16'h0B13;
		end
		32'h00006D8A: begin
				q			<=			16'hFFEB;
		end
		32'h00006D8C: begin
				q			<=			16'h0C13;
		end
		32'h00006D8E: begin
				q			<=			16'hFD50;
		end
		32'h00006D90: begin
				q			<=			16'h5783;
		end
		32'h00006D92: begin
				q			<=			16'h0D81;
		end
		32'h00006D94: begin
				q			<=			16'hF793;
		end
		32'h00006D96: begin
				q			<=			16'h0077;
		end
		32'h00006D98: begin
				q			<=			16'h9263;
		end
		32'h00006D9A: begin
				q			<=			16'h0607;
		end
		32'h00006D9C: begin
				q			<=			16'h0593;
		end
		32'h00006D9E: begin
				q			<=			16'h0A41;
		end
		32'h00006DA0: begin
				q			<=			16'h0513;
		end
		32'h00006DA2: begin
				q			<=			16'h0C01;
		end
		32'h00006DA4: begin
				q			<=			16'hE0EF;
		end
		32'h00006DA6: begin
				q			<=			16'hC98F;
		end
		32'h00006DA8: begin
				q			<=			16'h0513;
		end
		32'h00006DAA: begin
				q			<=			16'h0A41;
		end
		32'h00006DAC: begin
				q			<=			16'hE0EF;
		end
		32'h00006DAE: begin
				q			<=			16'hCF0F;
		end
		32'h00006DB0: begin
				q			<=			16'h0513;
		end
		32'h00006DB2: begin
				q			<=			16'h0A41;
		end
		32'h00006DB4: begin
				q			<=			16'hE0EF;
		end
		32'h00006DB6: begin
				q			<=			16'hCE8F;
		end
		32'h00006DB8: begin
				q			<=			16'h0593;
		end
		32'h00006DBA: begin
				q			<=			16'h0A41;
		end
		32'h00006DBC: begin
				q			<=			16'h0513;
		end
		32'h00006DBE: begin
				q			<=			16'h0C01;
		end
		32'h00006DC0: begin
				q			<=			16'hE0EF;
		end
		32'h00006DC2: begin
				q			<=			16'hE24F;
		end
		32'h00006DC4: begin
				q			<=			16'h5783;
		end
		32'h00006DC6: begin
				q			<=			16'h0A61;
		end
		32'h00006DC8: begin
				q			<=			16'h8793;
		end
		32'h00006DCA: begin
				q			<=			16'h0037;
		end
		32'h00006DCC: begin
				q			<=			16'h1323;
		end
		32'h00006DCE: begin
				q			<=			16'h0AF1;
		end
		32'h00006DD0: begin
				q			<=			16'h5783;
		end
		32'h00006DD2: begin
				q			<=			16'h0A81;
		end
		32'h00006DD4: begin
				q			<=			16'h9063;
		end
		32'h00006DD6: begin
				q			<=			16'h1207;
		end
		32'h00006DD8: begin
				q			<=			16'h5783;
		end
		32'h00006DDA: begin
				q			<=			16'h0BC1;
		end
		32'h00006DDC: begin
				q			<=			16'h9063;
		end
		32'h00006DDE: begin
				q			<=			16'h0207;
		end
		32'h00006DE0: begin
				q			<=			16'h5783;
		end
		32'h00006DE2: begin
				q			<=			16'h0A61;
		end
		32'h00006DE4: begin
				q			<=			16'h6C63;
		end
		32'h00006DE6: begin
				q			<=			16'h00FB;
		end
		32'h00006DE8: begin
				q			<=			16'h0593;
		end
		32'h00006DEA: begin
				q			<=			16'h0C01;
		end
		32'h00006DEC: begin
				q			<=			16'h0513;
		end
		32'h00006DEE: begin
				q			<=			16'h0A41;
		end
		32'h00006DF0: begin
				q			<=			16'h0413;
		end
		32'h00006DF2: begin
				q			<=			16'hFFF4;
		end
		32'h00006DF4: begin
				q			<=			16'hE0EF;
		end
		32'h00006DF6: begin
				q			<=			16'hC48F;
		end
		32'h00006DF8: begin
				q			<=			16'h1CE3;
		end
		32'h00006DFA: begin
				q			<=			16'hF984;
		end
		32'h00006DFC: begin
				q			<=			16'h0593;
		end
		32'h00006DFE: begin
				q			<=			16'h06C1;
		end
		32'h00006E00: begin
				q			<=			16'h0513;
		end
		32'h00006E02: begin
				q			<=			16'h0C01;
		end
		32'h00006E04: begin
				q			<=			16'hE0EF;
		end
		32'h00006E06: begin
				q			<=			16'hC0DF;
		end
		32'h00006E08: begin
				q			<=			16'h006F;
		end
		32'h00006E0A: begin
				q			<=			16'h0240;
		end
		32'h00006E0C: begin
				q			<=			16'h0613;
		end
		32'h00006E0E: begin
				q			<=			16'h06C1;
		end
		32'h00006E10: begin
				q			<=			16'h0693;
		end
		32'h00006E12: begin
				q			<=			16'h1501;
		end
		32'h00006E14: begin
				q			<=			16'h0593;
		end
		32'h00006E16: begin
				q			<=			16'h0006;
		end
		32'h00006E18: begin
				q			<=			16'h0513;
		end
		32'h00006E1A: begin
				q			<=			16'h000B;
		end
		32'h00006E1C: begin
				q			<=			16'hF0EF;
		end
		32'h00006E1E: begin
				q			<=			16'h99CF;
		end
		32'h00006E20: begin
				q			<=			16'h0413;
		end
		32'h00006E22: begin
				q			<=			16'hFFF4;
		end
		32'h00006E24: begin
				q			<=			16'h1783;
		end
		32'h00006E26: begin
				q			<=			16'h07C1;
		end
		32'h00006E28: begin
				q			<=			16'hD2E3;
		end
		32'h00006E2A: begin
				q			<=			16'hFE07;
		end
		32'h00006E2C: begin
				q			<=			16'h0593;
		end
		32'h00006E2E: begin
				q			<=			16'h0C01;
		end
		32'h00006E30: begin
				q			<=			16'h0513;
		end
		32'h00006E32: begin
				q			<=			16'h06C1;
		end
		32'h00006E34: begin
				q			<=			16'hE0EF;
		end
		32'h00006E36: begin
				q			<=			16'hBD8F;
		end
		32'h00006E38: begin
				q			<=			16'h0593;
		end
		32'h00006E3A: begin
				q			<=			16'h0881;
		end
		32'h00006E3C: begin
				q			<=			16'h8517;
		end
		32'h00006E3E: begin
				q			<=			16'h0000;
		end
		32'h00006E40: begin
				q			<=			16'h0513;
		end
		32'h00006E42: begin
				q			<=			16'h4845;
		end
		32'h00006E44: begin
				q			<=			16'hE0EF;
		end
		32'h00006E46: begin
				q			<=			16'hBC8F;
		end
		32'h00006E48: begin
				q			<=			16'h0C93;
		end
		32'h00006E4A: begin
				q			<=			16'h0000;
		end
		32'h00006E4C: begin
				q			<=			16'hFB37;
		end
		32'h00006E4E: begin
				q			<=			16'hFFFF;
		end
		32'h00006E50: begin
				q			<=			16'h0D13;
		end
		32'h00006E52: begin
				q			<=			16'h0020;
		end
		32'h00006E54: begin
				q			<=			16'h0D93;
		end
		32'h00006E56: begin
				q			<=			16'h1040;
		end
		32'h00006E58: begin
				q			<=			16'h8797;
		end
		32'h00006E5A: begin
				q			<=			16'h0000;
		end
		32'h00006E5C: begin
				q			<=			16'h8793;
		end
		32'h00006E5E: begin
				q			<=			16'h47C7;
		end
		32'h00006E60: begin
				q			<=			16'h8C33;
		end
		32'h00006E62: begin
				q			<=			16'h0197;
		end
		32'h00006E64: begin
				q			<=			16'h8797;
		end
		32'h00006E66: begin
				q			<=			16'h0000;
		end
		32'h00006E68: begin
				q			<=			16'h8793;
		end
		32'h00006E6A: begin
				q			<=			16'h5987;
		end
		32'h00006E6C: begin
				q			<=			16'h8733;
		end
		32'h00006E6E: begin
				q			<=			16'h0197;
		end
		32'h00006E70: begin
				q			<=			16'h0593;
		end
		32'h00006E72: begin
				q			<=			16'h0C01;
		end
		32'h00006E74: begin
				q			<=			16'h8517;
		end
		32'h00006E76: begin
				q			<=			16'h0000;
		end
		32'h00006E78: begin
				q			<=			16'h0513;
		end
		32'h00006E7A: begin
				q			<=			16'h44C5;
		end
		32'h00006E7C: begin
				q			<=			16'h2A23;
		end
		32'h00006E7E: begin
				q			<=			16'h00E1;
		end
		32'h00006E80: begin
				q			<=			16'hE0EF;
		end
		32'h00006E82: begin
				q			<=			16'hFB0F;
		end
		32'h00006E84: begin
				q			<=			16'h2703;
		end
		32'h00006E86: begin
				q			<=			16'h0141;
		end
		32'h00006E88: begin
				q			<=			16'h5663;
		end
		32'h00006E8A: begin
				q			<=			16'h04A0;
		end
		32'h00006E8C: begin
				q			<=			16'h0593;
		end
		32'h00006E8E: begin
				q			<=			16'h0C01;
		end
		32'h00006E90: begin
				q			<=			16'h0513;
		end
		32'h00006E92: begin
				q			<=			16'h0007;
		end
		32'h00006E94: begin
				q			<=			16'hE0EF;
		end
		32'h00006E96: begin
				q			<=			16'hF9CF;
		end
		32'h00006E98: begin
				q			<=			16'h4863;
		end
		32'h00006E9A: begin
				q			<=			16'h0205;
		end
		32'h00006E9C: begin
				q			<=			16'h0613;
		end
		32'h00006E9E: begin
				q			<=			16'h0C01;
		end
		32'h00006EA0: begin
				q			<=			16'h0593;
		end
		32'h00006EA2: begin
				q			<=			16'h0006;
		end
		32'h00006EA4: begin
				q			<=			16'h0693;
		end
		32'h00006EA6: begin
				q			<=			16'h1501;
		end
		32'h00006EA8: begin
				q			<=			16'h0513;
		end
		32'h00006EAA: begin
				q			<=			16'h000C;
		end
		32'h00006EAC: begin
				q			<=			16'hF0EF;
		end
		32'h00006EAE: begin
				q			<=			16'h90CF;
		end
		32'h00006EB0: begin
				q			<=			16'h0613;
		end
		32'h00006EB2: begin
				q			<=			16'h0881;
		end
		32'h00006EB4: begin
				q			<=			16'h0693;
		end
		32'h00006EB6: begin
				q			<=			16'h1501;
		end
		32'h00006EB8: begin
				q			<=			16'h0593;
		end
		32'h00006EBA: begin
				q			<=			16'h0006;
		end
		32'h00006EBC: begin
				q			<=			16'h0513;
		end
		32'h00006EBE: begin
				q			<=			16'h000C;
		end
		32'h00006EC0: begin
				q			<=			16'hF0EF;
		end
		32'h00006EC2: begin
				q			<=			16'h8F8F;
		end
		32'h00006EC4: begin
				q			<=			16'h0433;
		end
		32'h00006EC6: begin
				q			<=			16'h0164;
		end
		32'h00006EC8: begin
				q			<=			16'h8C93;
		end
		32'h00006ECA: begin
				q			<=			16'h014C;
		end
		32'h00006ECC: begin
				q			<=			16'h4B33;
		end
		32'h00006ECE: begin
				q			<=			16'h03AB;
		end
		32'h00006ED0: begin
				q			<=			16'h94E3;
		end
		32'h00006ED2: begin
				q			<=			16'hF9BC;
		end
		32'h00006ED4: begin
				q			<=			16'h0613;
		end
		32'h00006ED6: begin
				q			<=			16'h0881;
		end
		32'h00006ED8: begin
				q			<=			16'h0693;
		end
		32'h00006EDA: begin
				q			<=			16'h1501;
		end
		32'h00006EDC: begin
				q			<=			16'h8597;
		end
		32'h00006EDE: begin
				q			<=			16'h0000;
		end
		32'h00006EE0: begin
				q			<=			16'h8593;
		end
		32'h00006EE2: begin
				q			<=			16'h3E45;
		end
		32'h00006EE4: begin
				q			<=			16'h0513;
		end
		32'h00006EE6: begin
				q			<=			16'h0006;
		end
		32'h00006EE8: begin
				q			<=			16'hF097;
		end
		32'h00006EEA: begin
				q			<=			16'hFFFF;
		end
		32'h00006EEC: begin
				q			<=			16'h80E7;
		end
		32'h00006EEE: begin
				q			<=			16'h3AC0;
		end
		32'h00006EF0: begin
				q			<=			16'hF06F;
		end
		32'h00006EF2: begin
				q			<=			16'h8ADF;
		end
		32'h00006EF4: begin
				q			<=			16'h0513;
		end
		32'h00006EF6: begin
				q			<=			16'h0A41;
		end
		32'h00006EF8: begin
				q			<=			16'hE0EF;
		end
		32'h00006EFA: begin
				q			<=			16'hBA4F;
		end
		32'h00006EFC: begin
				q			<=			16'h5783;
		end
		32'h00006EFE: begin
				q			<=			16'h0A61;
		end
		32'h00006F00: begin
				q			<=			16'h8793;
		end
		32'h00006F02: begin
				q			<=			16'h0017;
		end
		32'h00006F04: begin
				q			<=			16'hF06F;
		end
		32'h00006F06: begin
				q			<=			16'hEC9F;
		end
		32'h00006F08: begin
				q			<=			16'h0513;
		end
		32'h00006F0A: begin
				q			<=			16'h06C1;
		end
		32'h00006F0C: begin
				q			<=			16'hE097;
		end
		32'h00006F0E: begin
				q			<=			16'hFFFF;
		end
		32'h00006F10: begin
				q			<=			16'h80E7;
		end
		32'h00006F12: begin
				q			<=			16'h3E00;
		end
		32'h00006F14: begin
				q			<=			16'h0593;
		end
		32'h00006F16: begin
				q			<=			16'h0A41;
		end
		32'h00006F18: begin
				q			<=			16'h0513;
		end
		32'h00006F1A: begin
				q			<=			16'h06C1;
		end
		32'h00006F1C: begin
				q			<=			16'hE0EF;
		end
		32'h00006F1E: begin
				q			<=			16'hB20F;
		end
		32'h00006F20: begin
				q			<=			16'h0513;
		end
		32'h00006F22: begin
				q			<=			16'h0A41;
		end
		32'h00006F24: begin
				q			<=			16'hE097;
		end
		32'h00006F26: begin
				q			<=			16'hFFFF;
		end
		32'h00006F28: begin
				q			<=			16'h80E7;
		end
		32'h00006F2A: begin
				q			<=			16'h3C80;
		end
		32'h00006F2C: begin
				q			<=			16'h0513;
		end
		32'h00006F2E: begin
				q			<=			16'h0A41;
		end
		32'h00006F30: begin
				q			<=			16'hE097;
		end
		32'h00006F32: begin
				q			<=			16'hFFFF;
		end
		32'h00006F34: begin
				q			<=			16'h80E7;
		end
		32'h00006F36: begin
				q			<=			16'h3BC0;
		end
		32'h00006F38: begin
				q			<=			16'h0593;
		end
		32'h00006F3A: begin
				q			<=			16'h06C1;
		end
		32'h00006F3C: begin
				q			<=			16'h0513;
		end
		32'h00006F3E: begin
				q			<=			16'h0A41;
		end
		32'h00006F40: begin
				q			<=			16'hE0EF;
		end
		32'h00006F42: begin
				q			<=			16'hCA4F;
		end
		32'h00006F44: begin
				q			<=			16'h0613;
		end
		32'h00006F46: begin
				q			<=			16'h1501;
		end
		32'h00006F48: begin
				q			<=			16'h0593;
		end
		32'h00006F4A: begin
				q			<=			16'h06C1;
		end
		32'h00006F4C: begin
				q			<=			16'h0513;
		end
		32'h00006F4E: begin
				q			<=			16'h0881;
		end
		32'h00006F50: begin
				q			<=			16'hF097;
		end
		32'h00006F52: begin
				q			<=			16'hFFFF;
		end
		32'h00006F54: begin
				q			<=			16'h80E7;
		end
		32'h00006F56: begin
				q			<=			16'hF780;
		end
		32'h00006F58: begin
				q			<=			16'h0413;
		end
		32'h00006F5A: begin
				q			<=			16'hFFF4;
		end
		32'h00006F5C: begin
				q			<=			16'h5B03;
		end
		32'h00006F5E: begin
				q			<=			16'h19C1;
		end
		32'h00006F60: begin
				q			<=			16'hF06F;
		end
		32'h00006F62: begin
				q			<=			16'h895F;
		end
		32'h00006F64: begin
				q			<=			16'h0B13;
		end
		32'h00006F66: begin
				q			<=			16'h030B;
		end
		32'h00006F68: begin
				q			<=			16'h0793;
		end
		32'h00006F6A: begin
				q			<=			16'h02E0;
		end
		32'h00006F6C: begin
				q			<=			16'h0AA3;
		end
		32'h00006F6E: begin
				q			<=			16'h1161;
		end
		32'h00006F70: begin
				q			<=			16'h0B23;
		end
		32'h00006F72: begin
				q			<=			16'h10F1;
		end
		32'h00006F74: begin
				q			<=			16'h0B13;
		end
		32'h00006F76: begin
				q			<=			16'h1171;
		end
		32'h00006F78: begin
				q			<=			16'h0A93;
		end
		32'h00006F7A: begin
				q			<=			16'h000B;
		end
		32'h00006F7C: begin
				q			<=			16'h87B3;
		end
		32'h00006F7E: begin
				q			<=			16'h416A;
		end
		32'h00006F80: begin
				q			<=			16'h5663;
		end
		32'h00006F82: begin
				q			<=			16'h04FC;
		end
		32'h00006F84: begin
				q			<=			16'h5783;
		end
		32'h00006F86: begin
				q			<=			16'h19C1;
		end
		32'h00006F88: begin
				q			<=			16'h0713;
		end
		32'h00006F8A: begin
				q			<=			16'h0040;
		end
		32'h00006F8C: begin
				q			<=			16'h8B13;
		end
		32'h00006F8E: begin
				q			<=			16'hFFFA;
		end
		32'h00006F90: begin
				q			<=			16'h5CE3;
		end
		32'h00006F92: begin
				q			<=			16'h8CF7;
		end
		32'h00006F94: begin
				q			<=			16'h0713;
		end
		32'h00006F96: begin
				q			<=			16'h0050;
		end
		32'h00006F98: begin
				q			<=			16'h8C63;
		end
		32'h00006F9A: begin
				q			<=			16'h08E7;
		end
		32'h00006F9C: begin
				q			<=			16'h0793;
		end
		32'h00006F9E: begin
				q			<=			16'h000B;
		end
		32'h00006FA0: begin
				q			<=			16'h0613;
		end
		32'h00006FA2: begin
				q			<=			16'h02E0;
		end
		32'h00006FA4: begin
				q			<=			16'h0593;
		end
		32'h00006FA6: begin
				q			<=			16'h0380;
		end
		32'h00006FA8: begin
				q			<=			16'h0693;
		end
		32'h00006FAA: begin
				q			<=			16'h0300;
		end
		32'h00006FAC: begin
				q			<=			16'h8793;
		end
		32'h00006FAE: begin
				q			<=			16'hFFF7;
		end
		32'h00006FB0: begin
				q			<=			16'hC703;
		end
		32'h00006FB2: begin
				q			<=			16'h0007;
		end
		32'h00006FB4: begin
				q			<=			16'h7713;
		end
		32'h00006FB6: begin
				q			<=			16'h07F7;
		end
		32'h00006FB8: begin
				q			<=			16'h5063;
		end
		32'h00006FBA: begin
				q			<=			16'h0C0C;
		end
		32'h00006FBC: begin
				q			<=			16'h0713;
		end
		32'h00006FBE: begin
				q			<=			16'h0310;
		end
		32'h00006FC0: begin
				q			<=			16'h8023;
		end
		32'h00006FC2: begin
				q			<=			16'h00E7;
		end
		32'h00006FC4: begin
				q			<=			16'h0413;
		end
		32'h00006FC6: begin
				q			<=			16'h0014;
		end
		32'h00006FC8: begin
				q			<=			16'hF06F;
		end
		32'h00006FCA: begin
				q			<=			16'h8A1F;
		end
		32'h00006FCC: begin
				q			<=			16'h0513;
		end
		32'h00006FCE: begin
				q			<=			16'h06C1;
		end
		32'h00006FD0: begin
				q			<=			16'hE097;
		end
		32'h00006FD2: begin
				q			<=			16'hFFFF;
		end
		32'h00006FD4: begin
				q			<=			16'h80E7;
		end
		32'h00006FD6: begin
				q			<=			16'h31C0;
		end
		32'h00006FD8: begin
				q			<=			16'h0593;
		end
		32'h00006FDA: begin
				q			<=			16'h0A41;
		end
		32'h00006FDC: begin
				q			<=			16'h0513;
		end
		32'h00006FDE: begin
				q			<=			16'h06C1;
		end
		32'h00006FE0: begin
				q			<=			16'hE0EF;
		end
		32'h00006FE2: begin
				q			<=			16'hA5CF;
		end
		32'h00006FE4: begin
				q			<=			16'h0513;
		end
		32'h00006FE6: begin
				q			<=			16'h0A41;
		end
		32'h00006FE8: begin
				q			<=			16'hE097;
		end
		32'h00006FEA: begin
				q			<=			16'hFFFF;
		end
		32'h00006FEC: begin
				q			<=			16'h80E7;
		end
		32'h00006FEE: begin
				q			<=			16'h3040;
		end
		32'h00006FF0: begin
				q			<=			16'h0513;
		end
		32'h00006FF2: begin
				q			<=			16'h0A41;
		end
		32'h00006FF4: begin
				q			<=			16'hE097;
		end
		32'h00006FF6: begin
				q			<=			16'hFFFF;
		end
		32'h00006FF8: begin
				q			<=			16'h80E7;
		end
		32'h00006FFA: begin
				q			<=			16'h2F80;
		end
		32'h00006FFC: begin
				q			<=			16'h0593;
		end
		32'h00006FFE: begin
				q			<=			16'h06C1;
		end
		32'h00007000: begin
				q			<=			16'h0513;
		end
		32'h00007002: begin
				q			<=			16'h0A41;
		end
		32'h00007004: begin
				q			<=			16'hE0EF;
		end
		32'h00007006: begin
				q			<=			16'hBE0F;
		end
		32'h00007008: begin
				q			<=			16'h0613;
		end
		32'h0000700A: begin
				q			<=			16'h1501;
		end
		32'h0000700C: begin
				q			<=			16'h0593;
		end
		32'h0000700E: begin
				q			<=			16'h06C1;
		end
		32'h00007010: begin
				q			<=			16'h0513;
		end
		32'h00007012: begin
				q			<=			16'h0881;
		end
		32'h00007014: begin
				q			<=			16'hF097;
		end
		32'h00007016: begin
				q			<=			16'hFFFF;
		end
		32'h00007018: begin
				q			<=			16'h80E7;
		end
		32'h0000701A: begin
				q			<=			16'hEB40;
		end
		32'h0000701C: begin
				q			<=			16'h4783;
		end
		32'h0000701E: begin
				q			<=			16'h19C1;
		end
		32'h00007020: begin
				q			<=			16'h8A93;
		end
		32'h00007022: begin
				q			<=			16'h001A;
		end
		32'h00007024: begin
				q			<=			16'h8793;
		end
		32'h00007026: begin
				q			<=			16'h0307;
		end
		32'h00007028: begin
				q			<=			16'h8FA3;
		end
		32'h0000702A: begin
				q			<=			16'hFEFA;
		end
		32'h0000702C: begin
				q			<=			16'hF06F;
		end
		32'h0000702E: begin
				q			<=			16'hF51F;
		end
		32'h00007030: begin
				q			<=			16'h0593;
		end
		32'h00007032: begin
				q			<=			16'h0881;
		end
		32'h00007034: begin
				q			<=			16'h0513;
		end
		32'h00007036: begin
				q			<=			16'h06C1;
		end
		32'h00007038: begin
				q			<=			16'hE0EF;
		end
		32'h0000703A: begin
				q			<=			16'h9D9F;
		end
		32'h0000703C: begin
				q			<=			16'h8597;
		end
		32'h0000703E: begin
				q			<=			16'h0000;
		end
		32'h00007040: begin
				q			<=			16'h8593;
		end
		32'h00007042: begin
				q			<=			16'h2705;
		end
		32'h00007044: begin
				q			<=			16'h0513;
		end
		32'h00007046: begin
				q			<=			16'h0881;
		end
		32'h00007048: begin
				q			<=			16'hE0EF;
		end
		32'h0000704A: begin
				q			<=			16'hDE8F;
		end
		32'h0000704C: begin
				q			<=			16'h18E3;
		end
		32'h0000704E: begin
				q			<=			16'hF405;
		end
		32'h00007050: begin
				q			<=			16'h4CE3;
		end
		32'h00007052: begin
				q			<=			16'h800C;
		end
		32'h00007054: begin
				q			<=			16'hC783;
		end
		32'h00007056: begin
				q			<=			16'hFFEA;
		end
		32'h00007058: begin
				q			<=			16'h8793;
		end
		32'h0000705A: begin
				q			<=			16'hFD27;
		end
		32'h0000705C: begin
				q			<=			16'hB793;
		end
		32'h0000705E: begin
				q			<=			16'h0017;
		end
		32'h00007060: begin
				q			<=			16'hC793;
		end
		32'h00007062: begin
				q			<=			16'hFFF7;
		end
		32'h00007064: begin
				q			<=			16'h07B3;
		end
		32'h00007066: begin
				q			<=			16'h00FB;
		end
		32'h00007068: begin
				q			<=			16'hC783;
		end
		32'h0000706A: begin
				q			<=			16'h0007;
		end
		32'h0000706C: begin
				q			<=			16'hF793;
		end
		32'h0000706E: begin
				q			<=			16'h0017;
		end
		32'h00007070: begin
				q			<=			16'h8C63;
		end
		32'h00007072: begin
				q			<=			16'hFE07;
		end
		32'h00007074: begin
				q			<=			16'hF06F;
		end
		32'h00007076: begin
				q			<=			16'hF29F;
		end
		32'h00007078: begin
				q			<=			16'h1463;
		end
		32'h0000707A: begin
				q			<=			16'h02C7;
		end
		32'h0000707C: begin
				q			<=			16'hC703;
		end
		32'h0000707E: begin
				q			<=			16'hFFF7;
		end
		32'h00007080: begin
				q			<=			16'h0693;
		end
		32'h00007082: begin
				q			<=			16'h0380;
		end
		32'h00007084: begin
				q			<=			16'hE863;
		end
		32'h00007086: begin
				q			<=			16'h00E6;
		end
		32'h00007088: begin
				q			<=			16'h0713;
		end
		32'h0000708A: begin
				q			<=			16'h0017;
		end
		32'h0000708C: begin
				q			<=			16'h8FA3;
		end
		32'h0000708E: begin
				q			<=			16'hFEE7;
		end
		32'h00007090: begin
				q			<=			16'hF06F;
		end
		32'h00007092: begin
				q			<=			16'hFD8F;
		end
		32'h00007094: begin
				q			<=			16'h0413;
		end
		32'h00007096: begin
				q			<=			16'h0014;
		end
		32'h00007098: begin
				q			<=			16'h0713;
		end
		32'h0000709A: begin
				q			<=			16'h0310;
		end
		32'h0000709C: begin
				q			<=			16'hF06F;
		end
		32'h0000709E: begin
				q			<=			16'hFF1F;
		end
		32'h000070A0: begin
				q			<=			16'hE863;
		end
		32'h000070A2: begin
				q			<=			16'h00E5;
		end
		32'h000070A4: begin
				q			<=			16'h0713;
		end
		32'h000070A6: begin
				q			<=			16'h0017;
		end
		32'h000070A8: begin
				q			<=			16'h8023;
		end
		32'h000070AA: begin
				q			<=			16'h00E7;
		end
		32'h000070AC: begin
				q			<=			16'hF06F;
		end
		32'h000070AE: begin
				q			<=			16'hFBCF;
		end
		32'h000070B0: begin
				q			<=			16'h8023;
		end
		32'h000070B2: begin
				q			<=			16'h00D7;
		end
		32'h000070B4: begin
				q			<=			16'hF06F;
		end
		32'h000070B6: begin
				q			<=			16'hEF9F;
		end
		32'h000070B8: begin
				q			<=			16'h0413;
		end
		32'h000070BA: begin
				q			<=			16'h0014;
		end
		32'h000070BC: begin
				q			<=			16'hA023;
		end
		32'h000070BE: begin
				q			<=			16'h008B;
		end
		32'h000070C0: begin
				q			<=			16'h8793;
		end
		32'h000070C2: begin
				q			<=			16'h000A;
		end
		32'h000070C4: begin
				q			<=			16'h0693;
		end
		32'h000070C6: begin
				q			<=			16'h02E0;
		end
		32'h000070C8: begin
				q			<=			16'hC703;
		end
		32'h000070CA: begin
				q			<=			16'h0007;
		end
		32'h000070CC: begin
				q			<=			16'h1E63;
		end
		32'h000070CE: begin
				q			<=			16'h0007;
		end
		32'h000070D0: begin
				q			<=			16'h0713;
		end
		32'h000070D2: begin
				q			<=			16'h0450;
		end
		32'h000070D4: begin
				q			<=			16'hC683;
		end
		32'h000070D6: begin
				q			<=			16'h0007;
		end
		32'h000070D8: begin
				q			<=			16'h8463;
		end
		32'h000070DA: begin
				q			<=			16'h00E6;
		end
		32'h000070DC: begin
				q			<=			16'hE863;
		end
		32'h000070DE: begin
				q			<=			16'h02FA;
		end
		32'h000070E0: begin
				q			<=			16'h8023;
		end
		32'h000070E2: begin
				q			<=			16'h0007;
		end
		32'h000070E4: begin
				q			<=			16'h006F;
		end
		32'h000070E6: begin
				q			<=			16'h0C80;
		end
		32'h000070E8: begin
				q			<=			16'h0C63;
		end
		32'h000070EA: begin
				q			<=			16'h00D7;
		end
		32'h000070EC: begin
				q			<=			16'h8793;
		end
		32'h000070EE: begin
				q			<=			16'h0017;
		end
		32'h000070F0: begin
				q			<=			16'hF06F;
		end
		32'h000070F2: begin
				q			<=			16'hFD9F;
		end
		32'h000070F4: begin
				q			<=			16'hC703;
		end
		32'h000070F6: begin
				q			<=			16'h0017;
		end
		32'h000070F8: begin
				q			<=			16'h8793;
		end
		32'h000070FA: begin
				q			<=			16'h0017;
		end
		32'h000070FC: begin
				q			<=			16'h8FA3;
		end
		32'h000070FE: begin
				q			<=			16'hFEE7;
		end
		32'h00007100: begin
				q			<=			16'hC703;
		end
		32'h00007102: begin
				q			<=			16'h0007;
		end
		32'h00007104: begin
				q			<=			16'h18E3;
		end
		32'h00007106: begin
				q			<=			16'hFE07;
		end
		32'h00007108: begin
				q			<=			16'hF06F;
		end
		32'h0000710A: begin
				q			<=			16'hFC9F;
		end
		32'h0000710C: begin
				q			<=			16'h8793;
		end
		32'h0000710E: begin
				q			<=			16'hFFF7;
		end
		32'h00007110: begin
				q			<=			16'hF06F;
		end
		32'h00007112: begin
				q			<=			16'hFC5F;
		end
		32'h00007114: begin
				q			<=			16'h8793;
		end
		32'h00007116: begin
				q			<=			16'h0017;
		end
		32'h00007118: begin
				q			<=			16'h006F;
		end
		32'h0000711A: begin
				q			<=			16'h0A00;
		end
		32'h0000711C: begin
				q			<=			16'h8413;
		end
		32'h0000711E: begin
				q			<=			16'h0006;
		end
		32'h00007120: begin
				q			<=			16'h006F;
		end
		32'h00007122: begin
				q			<=			16'h0A80;
		end
		32'h00007124: begin
				q			<=			16'h0413;
		end
		32'h00007126: begin
				q			<=			16'hFFF4;
		end
		32'h00007128: begin
				q			<=			16'h0023;
		end
		32'h0000712A: begin
				q			<=			16'h0004;
		end
		32'h0000712C: begin
				q			<=			16'h006F;
		end
		32'h0000712E: begin
				q			<=			16'h0CC0;
		end
		32'h00007130: begin
				q			<=			16'h8593;
		end
		32'h00007132: begin
				q			<=			16'h0015;
		end
		32'h00007134: begin
				q			<=			16'h2223;
		end
		32'h00007136: begin
				q			<=			16'h04B9;
		end
		32'h00007138: begin
				q			<=			16'h9793;
		end
		32'h0000713A: begin
				q			<=			16'h0017;
		end
		32'h0000713C: begin
				q			<=			16'h006F;
		end
		32'h0000713E: begin
				q			<=			16'h1040;
		end
		32'h00007140: begin
				q			<=			16'h87B7;
		end
		32'h00007142: begin
				q			<=			16'h0000;
		end
		32'h00007144: begin
				q			<=			16'h8793;
		end
		32'h00007146: begin
				q			<=			16'hFFF7;
		end
		32'h00007148: begin
				q			<=			16'h1463;
		end
		32'h0000714A: begin
				q			<=			16'hF4F7;
		end
		32'h0000714C: begin
				q			<=			16'h9597;
		end
		32'h0000714E: begin
				q			<=			16'h0000;
		end
		32'h00007150: begin
				q			<=			16'h8593;
		end
		32'h00007152: begin
				q			<=			16'hC785;
		end
		32'h00007154: begin
				q			<=			16'h8663;
		end
		32'h00007156: begin
				q			<=			16'h000A;
		end
		32'h00007158: begin
				q			<=			16'h9597;
		end
		32'h0000715A: begin
				q			<=			16'h0000;
		end
		32'h0000715C: begin
				q			<=			16'h8593;
		end
		32'h0000715E: begin
				q			<=			16'hC605;
		end
		32'h00007160: begin
				q			<=			16'h0513;
		end
		32'h00007162: begin
				q			<=			16'h1141;
		end
		32'h00007164: begin
				q			<=			16'h2437;
		end
		32'h00007166: begin
				q			<=			16'h0000;
		end
		32'h00007168: begin
				q			<=			16'h10EF;
		end
		32'h0000716A: begin
				q			<=			16'h1550;
		end
		32'h0000716C: begin
				q			<=			16'h0413;
		end
		32'h0000716E: begin
				q			<=			16'h70F4;
		end
		32'h00007170: begin
				q			<=			16'h2783;
		end
		32'h00007172: begin
				q			<=			16'h0101;
		end
		32'h00007174: begin
				q			<=			16'h0513;
		end
		32'h00007176: begin
				q			<=			16'h0501;
		end
		32'h00007178: begin
				q			<=			16'h2023;
		end
		32'h0000717A: begin
				q			<=			16'h1681;
		end
		32'h0000717C: begin
				q			<=			16'h2A23;
		end
		32'h0000717E: begin
				q			<=			16'h14F1;
		end
		32'h00007180: begin
				q			<=			16'hE097;
		end
		32'h00007182: begin
				q			<=			16'hFFFF;
		end
		32'h00007184: begin
				q			<=			16'h80E7;
		end
		32'h00007186: begin
				q			<=			16'h5C80;
		end
		32'h00007188: begin
				q			<=			16'h0A93;
		end
		32'h0000718A: begin
				q			<=			16'h1141;
		end
		32'h0000718C: begin
				q			<=			16'h1A63;
		end
		32'h0000718E: begin
				q			<=			16'h0005;
		end
		32'h00007190: begin
				q			<=			16'h0513;
		end
		32'h00007192: begin
				q			<=			16'h0501;
		end
		32'h00007194: begin
				q			<=			16'hE097;
		end
		32'h00007196: begin
				q			<=			16'hFFFF;
		end
		32'h00007198: begin
				q			<=			16'h80E7;
		end
		32'h0000719A: begin
				q			<=			16'h35C0;
		end
		32'h0000719C: begin
				q			<=			16'h0EE3;
		end
		32'h0000719E: begin
				q			<=			16'hF005;
		end
		32'h000071A0: begin
				q			<=			16'h27B7;
		end
		32'h000071A2: begin
				q			<=			16'h0000;
		end
		32'h000071A4: begin
				q			<=			16'h8793;
		end
		32'h000071A6: begin
				q			<=			16'h70F7;
		end
		32'h000071A8: begin
				q			<=			16'hA023;
		end
		32'h000071AA: begin
				q			<=			16'h00FB;
		end
		32'h000071AC: begin
				q			<=			16'h8793;
		end
		32'h000071AE: begin
				q			<=			16'h000A;
		end
		32'h000071B0: begin
				q			<=			16'h0613;
		end
		32'h000071B2: begin
				q			<=			16'h0200;
		end
		32'h000071B4: begin
				q			<=			16'h0693;
		end
		32'h000071B6: begin
				q			<=			16'h02D0;
		end
		32'h000071B8: begin
				q			<=			16'hC703;
		end
		32'h000071BA: begin
				q			<=			16'h0007;
		end
		32'h000071BC: begin
				q			<=			16'h0CE3;
		end
		32'h000071BE: begin
				q			<=			16'hF4C7;
		end
		32'h000071C0: begin
				q			<=			16'h0AE3;
		end
		32'h000071C2: begin
				q			<=			16'hF4D7;
		end
		32'h000071C4: begin
				q			<=			16'h8413;
		end
		32'h000071C6: begin
				q			<=			16'h000A;
		end
		32'h000071C8: begin
				q			<=			16'h8793;
		end
		32'h000071CA: begin
				q			<=			16'h0017;
		end
		32'h000071CC: begin
				q			<=			16'hC703;
		end
		32'h000071CE: begin
				q			<=			16'hFFF7;
		end
		32'h000071D0: begin
				q			<=			16'h0693;
		end
		32'h000071D2: begin
				q			<=			16'h0014;
		end
		32'h000071D4: begin
				q			<=			16'h8FA3;
		end
		32'h000071D6: begin
				q			<=			16'hFEE6;
		end
		32'h000071D8: begin
				q			<=			16'h12E3;
		end
		32'h000071DA: begin
				q			<=			16'hF407;
		end
		32'h000071DC: begin
				q			<=			16'h0713;
		end
		32'h000071DE: begin
				q			<=			16'h0020;
		end
		32'h000071E0: begin
				q			<=			16'h0793;
		end
		32'h000071E2: begin
				q			<=			16'h0010;
		end
		32'h000071E4: begin
				q			<=			16'h0863;
		end
		32'h000071E6: begin
				q			<=			16'h00EA;
		end
		32'h000071E8: begin
				q			<=			16'h2783;
		end
		32'h000071EA: begin
				q			<=			16'h1601;
		end
		32'h000071EC: begin
				q			<=			16'hD463;
		end
		32'h000071EE: begin
				q			<=			16'h0097;
		end
		32'h000071F0: begin
				q			<=			16'h8793;
		end
		32'h000071F2: begin
				q			<=			16'h0004;
		end
		32'h000071F4: begin
				q			<=			16'h0693;
		end
		32'h000071F6: begin
				q			<=			16'h0300;
		end
		32'h000071F8: begin
				q			<=			16'h4703;
		end
		32'h000071FA: begin
				q			<=			16'hFFF4;
		end
		32'h000071FC: begin
				q			<=			16'h1663;
		end
		32'h000071FE: begin
				q			<=			16'h00D7;
		end
		32'h00007200: begin
				q			<=			16'h0733;
		end
		32'h00007202: begin
				q			<=			16'h4154;
		end
		32'h00007204: begin
				q			<=			16'hC0E3;
		end
		32'h00007206: begin
				q			<=			16'hF2E7;
		end
		32'h00007208: begin
				q			<=			16'h0793;
		end
		32'h0000720A: begin
				q			<=			16'h0030;
		end
		32'h0000720C: begin
				q			<=			16'h8713;
		end
		32'h0000720E: begin
				q			<=			16'h0099;
		end
		32'h00007210: begin
				q			<=			16'h1463;
		end
		32'h00007212: begin
				q			<=			16'h02FA;
		end
		32'h00007214: begin
				q			<=			16'h2783;
		end
		32'h00007216: begin
				q			<=			16'h1601;
		end
		32'h00007218: begin
				q			<=			16'h84B3;
		end
		32'h0000721A: begin
				q			<=			16'h00F4;
		end
		32'h0000721C: begin
				q			<=			16'hD863;
		end
		32'h0000721E: begin
				q			<=			16'h0004;
		end
		32'h00007220: begin
				q			<=			16'h0A23;
		end
		32'h00007222: begin
				q			<=			16'h1001;
		end
		32'h00007224: begin
				q			<=			16'hA023;
		end
		32'h00007226: begin
				q			<=			16'h000B;
		end
		32'h00007228: begin
				q			<=			16'h8413;
		end
		32'h0000722A: begin
				q			<=			16'h000A;
		end
		32'h0000722C: begin
				q			<=			16'hA783;
		end
		32'h0000722E: begin
				q			<=			16'h000B;
		end
		32'h00007230: begin
				q			<=			16'h89B3;
		end
		32'h00007232: begin
				q			<=			16'h00F9;
		end
		32'h00007234: begin
				q			<=			16'h8713;
		end
		32'h00007236: begin
				q			<=			16'h0039;
		end
		32'h00007238: begin
				q			<=			16'h2223;
		end
		32'h0000723A: begin
				q			<=			16'h0409;
		end
		32'h0000723C: begin
				q			<=			16'h0793;
		end
		32'h0000723E: begin
				q			<=			16'h0040;
		end
		32'h00007240: begin
				q			<=			16'h8693;
		end
		32'h00007242: begin
				q			<=			16'h0147;
		end
		32'h00007244: begin
				q			<=			16'h2583;
		end
		32'h00007246: begin
				q			<=			16'h0449;
		end
		32'h00007248: begin
				q			<=			16'h74E3;
		end
		32'h0000724A: begin
				q			<=			16'hEED7;
		end
		32'h0000724C: begin
				q			<=			16'h0513;
		end
		32'h0000724E: begin
				q			<=			16'h0009;
		end
		32'h00007250: begin
				q			<=			16'h1097;
		end
		32'h00007252: begin
				q			<=			16'h0000;
		end
		32'h00007254: begin
				q			<=			16'h80E7;
		end
		32'h00007256: begin
				q			<=			16'h83C0;
		end
		32'h00007258: begin
				q			<=			16'h2023;
		end
		32'h0000725A: begin
				q			<=			16'h04A9;
		end
		32'h0000725C: begin
				q			<=			16'h8593;
		end
		32'h0000725E: begin
				q			<=			16'h000A;
		end
		32'h00007260: begin
				q			<=			16'h0493;
		end
		32'h00007262: begin
				q			<=			16'h0005;
		end
		32'h00007264: begin
				q			<=			16'h2097;
		end
		32'h00007266: begin
				q			<=			16'h0000;
		end
		32'h00007268: begin
				q			<=			16'h80E7;
		end
		32'h0000726A: begin
				q			<=			16'h8D80;
		end
		32'h0000726C: begin
				q			<=			16'h2783;
		end
		32'h0000726E: begin
				q			<=			16'h00C1;
		end
		32'h00007270: begin
				q			<=			16'h8863;
		end
		32'h00007272: begin
				q			<=			16'h0007;
		end
		32'h00007274: begin
				q			<=			16'h0433;
		end
		32'h00007276: begin
				q			<=			16'h4154;
		end
		32'h00007278: begin
				q			<=			16'h8433;
		end
		32'h0000727A: begin
				q			<=			16'h0084;
		end
		32'h0000727C: begin
				q			<=			16'hA023;
		end
		32'h0000727E: begin
				q			<=			16'h0087;
		end
		32'h00007280: begin
				q			<=			16'h2083;
		end
		32'h00007282: begin
				q			<=			16'h1DC1;
		end
		32'h00007284: begin
				q			<=			16'h2403;
		end
		32'h00007286: begin
				q			<=			16'h1D81;
		end
		32'h00007288: begin
				q			<=			16'h8513;
		end
		32'h0000728A: begin
				q			<=			16'h0004;
		end
		32'h0000728C: begin
				q			<=			16'h2903;
		end
		32'h0000728E: begin
				q			<=			16'h1D01;
		end
		32'h00007290: begin
				q			<=			16'h2483;
		end
		32'h00007292: begin
				q			<=			16'h1D41;
		end
		32'h00007294: begin
				q			<=			16'h2983;
		end
		32'h00007296: begin
				q			<=			16'h1CC1;
		end
		32'h00007298: begin
				q			<=			16'h2A03;
		end
		32'h0000729A: begin
				q			<=			16'h1C81;
		end
		32'h0000729C: begin
				q			<=			16'h2A83;
		end
		32'h0000729E: begin
				q			<=			16'h1C41;
		end
		32'h000072A0: begin
				q			<=			16'h2B03;
		end
		32'h000072A2: begin
				q			<=			16'h1C01;
		end
		32'h000072A4: begin
				q			<=			16'h2B83;
		end
		32'h000072A6: begin
				q			<=			16'h1BC1;
		end
		32'h000072A8: begin
				q			<=			16'h2C03;
		end
		32'h000072AA: begin
				q			<=			16'h1B81;
		end
		32'h000072AC: begin
				q			<=			16'h2C83;
		end
		32'h000072AE: begin
				q			<=			16'h1B41;
		end
		32'h000072B0: begin
				q			<=			16'h2D03;
		end
		32'h000072B2: begin
				q			<=			16'h1B01;
		end
		32'h000072B4: begin
				q			<=			16'h2D83;
		end
		32'h000072B6: begin
				q			<=			16'h1AC1;
		end
		32'h000072B8: begin
				q			<=			16'h0113;
		end
		32'h000072BA: begin
				q			<=			16'h1E01;
		end
		32'h000072BC: begin
				q			<=			16'h8067;
		end
		32'h000072BE: begin
				q			<=			16'h0000;
		end
		32'h000072C0: begin
				q			<=			16'h0793;
		end
		32'h000072C2: begin
				q			<=			16'h00A0;
		end
		32'h000072C4: begin
				q			<=			16'h0C13;
		end
		32'h000072C6: begin
				q			<=			16'h02A0;
		end
		32'h000072C8: begin
				q			<=			16'h1EE3;
		end
		32'h000072CA: begin
				q			<=			16'hC8FB;
		end
		32'h000072CC: begin
				q			<=			16'h0793;
		end
		32'h000072CE: begin
				q			<=			16'h0310;
		end
		32'h000072D0: begin
				q			<=			16'h0AA3;
		end
		32'h000072D2: begin
				q			<=			16'h10F1;
		end
		32'h000072D4: begin
				q			<=			16'h0793;
		end
		32'h000072D6: begin
				q			<=			16'h02E0;
		end
		32'h000072D8: begin
				q			<=			16'h0B23;
		end
		32'h000072DA: begin
				q			<=			16'h10F1;
		end
		32'h000072DC: begin
				q			<=			16'h0C13;
		end
		32'h000072DE: begin
				q			<=			16'h02A0;
		end
		32'h000072E0: begin
				q			<=			16'hF06F;
		end
		32'h000072E2: begin
				q			<=			16'hD70F;
		end
		32'h000072E4: begin
				q			<=			16'h2783;
		end
		32'h000072E6: begin
				q			<=			16'h0005;
		end
		32'h000072E8: begin
				q			<=			16'h0113;
		end
		32'h000072EA: begin
				q			<=			16'hFC01;
		end
		32'h000072EC: begin
				q			<=			16'h0593;
		end
		32'h000072EE: begin
				q			<=			16'h0141;
		end
		32'h000072F0: begin
				q			<=			16'h2023;
		end
		32'h000072F2: begin
				q			<=			16'h00F1;
		end
		32'h000072F4: begin
				q			<=			16'h2783;
		end
		32'h000072F6: begin
				q			<=			16'h0045;
		end
		32'h000072F8: begin
				q			<=			16'h2E23;
		end
		32'h000072FA: begin
				q			<=			16'h0211;
		end
		32'h000072FC: begin
				q			<=			16'h2223;
		end
		32'h000072FE: begin
				q			<=			16'h00F1;
		end
		32'h00007300: begin
				q			<=			16'h2783;
		end
		32'h00007302: begin
				q			<=			16'h0085;
		end
		32'h00007304: begin
				q			<=			16'h2423;
		end
		32'h00007306: begin
				q			<=			16'h00F1;
		end
		32'h00007308: begin
				q			<=			16'h2783;
		end
		32'h0000730A: begin
				q			<=			16'h00C5;
		end
		32'h0000730C: begin
				q			<=			16'h0513;
		end
		32'h0000730E: begin
				q			<=			16'h0001;
		end
		32'h00007310: begin
				q			<=			16'h2623;
		end
		32'h00007312: begin
				q			<=			16'h00F1;
		end
		32'h00007314: begin
				q			<=			16'hE0EF;
		end
		32'h00007316: begin
				q			<=			16'hF70F;
		end
		32'h00007318: begin
				q			<=			16'h5783;
		end
		32'h0000731A: begin
				q			<=			16'h0261;
		end
		32'h0000731C: begin
				q			<=			16'h0513;
		end
		32'h0000731E: begin
				q			<=			16'h0000;
		end
		32'h00007320: begin
				q			<=			16'hC793;
		end
		32'h00007322: begin
				q			<=			16'hFFF7;
		end
		32'h00007324: begin
				q			<=			16'h9713;
		end
		32'h00007326: begin
				q			<=			16'h0117;
		end
		32'h00007328: begin
				q			<=			16'h1A63;
		end
		32'h0000732A: begin
				q			<=			16'h0007;
		end
		32'h0000732C: begin
				q			<=			16'h0513;
		end
		32'h0000732E: begin
				q			<=			16'h0141;
		end
		32'h00007330: begin
				q			<=			16'hE0EF;
		end
		32'h00007332: begin
				q			<=			16'h9C0F;
		end
		32'h00007334: begin
				q			<=			16'h3513;
		end
		32'h00007336: begin
				q			<=			16'h0015;
		end
		32'h00007338: begin
				q			<=			16'h0513;
		end
		32'h0000733A: begin
				q			<=			16'h0015;
		end
		32'h0000733C: begin
				q			<=			16'h2083;
		end
		32'h0000733E: begin
				q			<=			16'h03C1;
		end
		32'h00007340: begin
				q			<=			16'h0113;
		end
		32'h00007342: begin
				q			<=			16'h0401;
		end
		32'h00007344: begin
				q			<=			16'h8067;
		end
		32'h00007346: begin
				q			<=			16'h0000;
		end
		32'h00007348: begin
				q			<=			16'h0000;
		end
		32'h0000734A: begin
				q			<=			16'h0000;
		end
		32'h0000734C: begin
				q			<=			16'h0513;
		end
		32'h0000734E: begin
				q			<=			16'h0F05;
		end
		32'h00007350: begin
				q			<=			16'h8067;
		end
		32'h00007352: begin
				q			<=			16'h0000;
		end
		32'h00007354: begin
				q			<=			16'h9797;
		end
		32'h00007356: begin
				q			<=			16'h0000;
		end
		32'h00007358: begin
				q			<=			16'h8793;
		end
		32'h0000735A: begin
				q			<=			16'h5847;
		end
		32'h0000735C: begin
				q			<=			16'hA783;
		end
		32'h0000735E: begin
				q			<=			16'h0007;
		end
		32'h00007360: begin
				q			<=			16'hA503;
		end
		32'h00007362: begin
				q			<=			16'h0347;
		end
		32'h00007364: begin
				q			<=			16'h1663;
		end
		32'h00007366: begin
				q			<=			16'h0005;
		end
		32'h00007368: begin
				q			<=			16'h9517;
		end
		32'h0000736A: begin
				q			<=			16'h0000;
		end
		32'h0000736C: begin
				q			<=			16'h0513;
		end
		32'h0000736E: begin
				q			<=			16'h4005;
		end
		32'h00007370: begin
				q			<=			16'h0513;
		end
		32'h00007372: begin
				q			<=			16'h0F05;
		end
		32'h00007374: begin
				q			<=			16'h8067;
		end
		32'h00007376: begin
				q			<=			16'h0000;
		end
		32'h00007378: begin
				q			<=			16'h9797;
		end
		32'h0000737A: begin
				q			<=			16'h0000;
		end
		32'h0000737C: begin
				q			<=			16'h8793;
		end
		32'h0000737E: begin
				q			<=			16'h5607;
		end
		32'h00007380: begin
				q			<=			16'hA783;
		end
		32'h00007382: begin
				q			<=			16'h0007;
		end
		32'h00007384: begin
				q			<=			16'hA503;
		end
		32'h00007386: begin
				q			<=			16'h0347;
		end
		32'h00007388: begin
				q			<=			16'h1663;
		end
		32'h0000738A: begin
				q			<=			16'h0005;
		end
		32'h0000738C: begin
				q			<=			16'h9517;
		end
		32'h0000738E: begin
				q			<=			16'h0000;
		end
		32'h00007390: begin
				q			<=			16'h0513;
		end
		32'h00007392: begin
				q			<=			16'h3DC5;
		end
		32'h00007394: begin
				q			<=			16'h0513;
		end
		32'h00007396: begin
				q			<=			16'h0F05;
		end
		32'h00007398: begin
				q			<=			16'h8067;
		end
		32'h0000739A: begin
				q			<=			16'h0000;
		end
		32'h0000739C: begin
				q			<=			16'h0000;
		end
		32'h0000739E: begin
				q			<=			16'h0000;
		end
		32'h000073A0: begin
				q			<=			16'h0113;
		end
		32'h000073A2: begin
				q			<=			16'hFD01;
		end
		32'h000073A4: begin
				q			<=			16'h2623;
		end
		32'h000073A6: begin
				q			<=			16'h0211;
		end
		32'h000073A8: begin
				q			<=			16'h2423;
		end
		32'h000073AA: begin
				q			<=			16'h0281;
		end
		32'h000073AC: begin
				q			<=			16'h2223;
		end
		32'h000073AE: begin
				q			<=			16'h0291;
		end
		32'h000073B0: begin
				q			<=			16'h2023;
		end
		32'h000073B2: begin
				q			<=			16'h0321;
		end
		32'h000073B4: begin
				q			<=			16'h2E23;
		end
		32'h000073B6: begin
				q			<=			16'h0131;
		end
		32'h000073B8: begin
				q			<=			16'h2C23;
		end
		32'h000073BA: begin
				q			<=			16'h0141;
		end
		32'h000073BC: begin
				q			<=			16'h2A23;
		end
		32'h000073BE: begin
				q			<=			16'h0151;
		end
		32'h000073C0: begin
				q			<=			16'h2823;
		end
		32'h000073C2: begin
				q			<=			16'h0161;
		end
		32'h000073C4: begin
				q			<=			16'h2623;
		end
		32'h000073C6: begin
				q			<=			16'h0171;
		end
		32'h000073C8: begin
				q			<=			16'h2423;
		end
		32'h000073CA: begin
				q			<=			16'h0181;
		end
		32'h000073CC: begin
				q			<=			16'h8793;
		end
		32'h000073CE: begin
				q			<=			16'h00B5;
		end
		32'h000073D0: begin
				q			<=			16'h0713;
		end
		32'h000073D2: begin
				q			<=			16'h0160;
		end
		32'h000073D4: begin
				q			<=			16'h7463;
		end
		32'h000073D6: begin
				q			<=			16'h04F7;
		end
		32'h000073D8: begin
				q			<=			16'hF493;
		end
		32'h000073DA: begin
				q			<=			16'hFF87;
		end
		32'h000073DC: begin
				q			<=			16'hD263;
		end
		32'h000073DE: begin
				q			<=			16'h0404;
		end
		32'h000073E0: begin
				q			<=			16'h0793;
		end
		32'h000073E2: begin
				q			<=			16'h00C0;
		end
		32'h000073E4: begin
				q			<=			16'h2023;
		end
		32'h000073E6: begin
				q			<=			16'h00F5;
		end
		32'h000073E8: begin
				q			<=			16'h0513;
		end
		32'h000073EA: begin
				q			<=			16'h0000;
		end
		32'h000073EC: begin
				q			<=			16'h2083;
		end
		32'h000073EE: begin
				q			<=			16'h02C1;
		end
		32'h000073F0: begin
				q			<=			16'h2403;
		end
		32'h000073F2: begin
				q			<=			16'h0281;
		end
		32'h000073F4: begin
				q			<=			16'h2483;
		end
		32'h000073F6: begin
				q			<=			16'h0241;
		end
		32'h000073F8: begin
				q			<=			16'h2903;
		end
		32'h000073FA: begin
				q			<=			16'h0201;
		end
		32'h000073FC: begin
				q			<=			16'h2983;
		end
		32'h000073FE: begin
				q			<=			16'h01C1;
		end
		32'h00007400: begin
				q			<=			16'h2A03;
		end
		32'h00007402: begin
				q			<=			16'h0181;
		end
		32'h00007404: begin
				q			<=			16'h2A83;
		end
		32'h00007406: begin
				q			<=			16'h0141;
		end
		32'h00007408: begin
				q			<=			16'h2B03;
		end
		32'h0000740A: begin
				q			<=			16'h0101;
		end
		32'h0000740C: begin
				q			<=			16'h2B83;
		end
		32'h0000740E: begin
				q			<=			16'h00C1;
		end
		32'h00007410: begin
				q			<=			16'h2C03;
		end
		32'h00007412: begin
				q			<=			16'h0081;
		end
		32'h00007414: begin
				q			<=			16'h0113;
		end
		32'h00007416: begin
				q			<=			16'h0301;
		end
		32'h00007418: begin
				q			<=			16'h8067;
		end
		32'h0000741A: begin
				q			<=			16'h0000;
		end
		32'h0000741C: begin
				q			<=			16'h0493;
		end
		32'h0000741E: begin
				q			<=			16'h0100;
		end
		32'h00007420: begin
				q			<=			16'hE0E3;
		end
		32'h00007422: begin
				q			<=			16'hFCB4;
		end
		32'h00007424: begin
				q			<=			16'h0913;
		end
		32'h00007426: begin
				q			<=			16'h0005;
		end
		32'h00007428: begin
				q			<=			16'h00EF;
		end
		32'h0000742A: begin
				q			<=			16'h6580;
		end
		32'h0000742C: begin
				q			<=			16'h0793;
		end
		32'h0000742E: begin
				q			<=			16'h1F70;
		end
		32'h00007430: begin
				q			<=			16'h9997;
		end
		32'h00007432: begin
				q			<=			16'h0000;
		end
		32'h00007434: begin
				q			<=			16'h8993;
		end
		32'h00007436: begin
				q			<=			16'hF309;
		end
		32'h00007438: begin
				q			<=			16'hEA63;
		end
		32'h0000743A: begin
				q			<=			16'h0497;
		end
		32'h0000743C: begin
				q			<=			16'h8713;
		end
		32'h0000743E: begin
				q			<=			16'h0084;
		end
		32'h00007440: begin
				q			<=			16'h8733;
		end
		32'h00007442: begin
				q			<=			16'h00E9;
		end
		32'h00007444: begin
				q			<=			16'h2403;
		end
		32'h00007446: begin
				q			<=			16'h0047;
		end
		32'h00007448: begin
				q			<=			16'h0693;
		end
		32'h0000744A: begin
				q			<=			16'hFF87;
		end
		32'h0000744C: begin
				q			<=			16'hD793;
		end
		32'h0000744E: begin
				q			<=			16'h0034;
		end
		32'h00007450: begin
				q			<=			16'h1863;
		end
		32'h00007452: begin
				q			<=			16'h00D4;
		end
		32'h00007454: begin
				q			<=			16'h2403;
		end
		32'h00007456: begin
				q			<=			16'h00C7;
		end
		32'h00007458: begin
				q			<=			16'h8793;
		end
		32'h0000745A: begin
				q			<=			16'h0027;
		end
		32'h0000745C: begin
				q			<=			16'h0063;
		end
		32'h0000745E: begin
				q			<=			16'h0887;
		end
		32'h00007460: begin
				q			<=			16'h2783;
		end
		32'h00007462: begin
				q			<=			16'h0044;
		end
		32'h00007464: begin
				q			<=			16'h2703;
		end
		32'h00007466: begin
				q			<=			16'h00C4;
		end
		32'h00007468: begin
				q			<=			16'h2683;
		end
		32'h0000746A: begin
				q			<=			16'h0084;
		end
		32'h0000746C: begin
				q			<=			16'hF793;
		end
		32'h0000746E: begin
				q			<=			16'hFFC7;
		end
		32'h00007470: begin
				q			<=			16'h07B3;
		end
		32'h00007472: begin
				q			<=			16'h00F4;
		end
		32'h00007474: begin
				q			<=			16'hA623;
		end
		32'h00007476: begin
				q			<=			16'h00E6;
		end
		32'h00007478: begin
				q			<=			16'h2423;
		end
		32'h0000747A: begin
				q			<=			16'h00D7;
		end
		32'h0000747C: begin
				q			<=			16'hA703;
		end
		32'h0000747E: begin
				q			<=			16'h0047;
		end
		32'h00007480: begin
				q			<=			16'h6713;
		end
		32'h00007482: begin
				q			<=			16'h0017;
		end
		32'h00007484: begin
				q			<=			16'hA223;
		end
		32'h00007486: begin
				q			<=			16'h00E7;
		end
		32'h00007488: begin
				q			<=			16'h006F;
		end
		32'h0000748A: begin
				q			<=			16'h0AC0;
		end
		32'h0000748C: begin
				q			<=			16'hD713;
		end
		32'h0000748E: begin
				q			<=			16'h0094;
		end
		32'h00007490: begin
				q			<=			16'h0793;
		end
		32'h00007492: begin
				q			<=			16'h03F0;
		end
		32'h00007494: begin
				q			<=			16'h0A63;
		end
		32'h00007496: begin
				q			<=			16'h0007;
		end
		32'h00007498: begin
				q			<=			16'h0793;
		end
		32'h0000749A: begin
				q			<=			16'h0040;
		end
		32'h0000749C: begin
				q			<=			16'hE663;
		end
		32'h0000749E: begin
				q			<=			16'h0AE7;
		end
		32'h000074A0: begin
				q			<=			16'hD793;
		end
		32'h000074A2: begin
				q			<=			16'h0064;
		end
		32'h000074A4: begin
				q			<=			16'h8793;
		end
		32'h000074A6: begin
				q			<=			16'h0387;
		end
		32'h000074A8: begin
				q			<=			16'h8713;
		end
		32'h000074AA: begin
				q			<=			16'h0017;
		end
		32'h000074AC: begin
				q			<=			16'h1713;
		end
		32'h000074AE: begin
				q			<=			16'h0037;
		end
		32'h000074B0: begin
				q			<=			16'h8733;
		end
		32'h000074B2: begin
				q			<=			16'h00E9;
		end
		32'h000074B4: begin
				q			<=			16'h2403;
		end
		32'h000074B6: begin
				q			<=			16'h0047;
		end
		32'h000074B8: begin
				q			<=			16'h0593;
		end
		32'h000074BA: begin
				q			<=			16'hFF87;
		end
		32'h000074BC: begin
				q			<=			16'h0513;
		end
		32'h000074BE: begin
				q			<=			16'h00F0;
		end
		32'h000074C0: begin
				q			<=			16'h0C63;
		end
		32'h000074C2: begin
				q			<=			16'h00B4;
		end
		32'h000074C4: begin
				q			<=			16'h2703;
		end
		32'h000074C6: begin
				q			<=			16'h0044;
		end
		32'h000074C8: begin
				q			<=			16'h7713;
		end
		32'h000074CA: begin
				q			<=			16'hFFC7;
		end
		32'h000074CC: begin
				q			<=			16'h0633;
		end
		32'h000074CE: begin
				q			<=			16'h4097;
		end
		32'h000074D0: begin
				q			<=			16'h5463;
		end
		32'h000074D2: begin
				q			<=			16'h0CC5;
		end
		32'h000074D4: begin
				q			<=			16'h8793;
		end
		32'h000074D6: begin
				q			<=			16'hFFF7;
		end
		32'h000074D8: begin
				q			<=			16'h8793;
		end
		32'h000074DA: begin
				q			<=			16'h0017;
		end
		32'h000074DC: begin
				q			<=			16'hA403;
		end
		32'h000074DE: begin
				q			<=			16'h0109;
		end
		32'h000074E0: begin
				q			<=			16'h9597;
		end
		32'h000074E2: begin
				q			<=			16'h0000;
		end
		32'h000074E4: begin
				q			<=			16'h8593;
		end
		32'h000074E6: begin
				q			<=			16'hE885;
		end
		32'h000074E8: begin
				q			<=			16'h0463;
		end
		32'h000074EA: begin
				q			<=			16'h14B4;
		end
		32'h000074EC: begin
				q			<=			16'h2703;
		end
		32'h000074EE: begin
				q			<=			16'h0044;
		end
		32'h000074F0: begin
				q			<=			16'h0693;
		end
		32'h000074F2: begin
				q			<=			16'h00F0;
		end
		32'h000074F4: begin
				q			<=			16'h7713;
		end
		32'h000074F6: begin
				q			<=			16'hFFC7;
		end
		32'h000074F8: begin
				q			<=			16'h0633;
		end
		32'h000074FA: begin
				q			<=			16'h4097;
		end
		32'h000074FC: begin
				q			<=			16'hD063;
		end
		32'h000074FE: begin
				q			<=			16'h0CC6;
		end
		32'h00007500: begin
				q			<=			16'hE793;
		end
		32'h00007502: begin
				q			<=			16'h0014;
		end
		32'h00007504: begin
				q			<=			16'h2223;
		end
		32'h00007506: begin
				q			<=			16'h00F4;
		end
		32'h00007508: begin
				q			<=			16'h06B3;
		end
		32'h0000750A: begin
				q			<=			16'h0094;
		end
		32'h0000750C: begin
				q			<=			16'h9797;
		end
		32'h0000750E: begin
				q			<=			16'h0000;
		end
		32'h00007510: begin
				q			<=			16'hA423;
		end
		32'h00007512: begin
				q			<=			16'hE6D7;
		end
		32'h00007514: begin
				q			<=			16'h9797;
		end
		32'h00007516: begin
				q			<=			16'h0000;
		end
		32'h00007518: begin
				q			<=			16'hAE23;
		end
		32'h0000751A: begin
				q			<=			16'hE4D7;
		end
		32'h0000751C: begin
				q			<=			16'h6793;
		end
		32'h0000751E: begin
				q			<=			16'h0016;
		end
		32'h00007520: begin
				q			<=			16'hA623;
		end
		32'h00007522: begin
				q			<=			16'h00B6;
		end
		32'h00007524: begin
				q			<=			16'hA423;
		end
		32'h00007526: begin
				q			<=			16'h00B6;
		end
		32'h00007528: begin
				q			<=			16'hA223;
		end
		32'h0000752A: begin
				q			<=			16'h00F6;
		end
		32'h0000752C: begin
				q			<=			16'h0733;
		end
		32'h0000752E: begin
				q			<=			16'h00E4;
		end
		32'h00007530: begin
				q			<=			16'h2023;
		end
		32'h00007532: begin
				q			<=			16'h00C7;
		end
		32'h00007534: begin
				q			<=			16'h0513;
		end
		32'h00007536: begin
				q			<=			16'h0009;
		end
		32'h00007538: begin
				q			<=			16'h0097;
		end
		32'h0000753A: begin
				q			<=			16'h0000;
		end
		32'h0000753C: begin
				q			<=			16'h80E7;
		end
		32'h0000753E: begin
				q			<=			16'h54C0;
		end
		32'h00007540: begin
				q			<=			16'h0513;
		end
		32'h00007542: begin
				q			<=			16'h0084;
		end
		32'h00007544: begin
				q			<=			16'hF06F;
		end
		32'h00007546: begin
				q			<=			16'hEA9F;
		end
		32'h00007548: begin
				q			<=			16'h0793;
		end
		32'h0000754A: begin
				q			<=			16'h0140;
		end
		32'h0000754C: begin
				q			<=			16'hE663;
		end
		32'h0000754E: begin
				q			<=			16'h00E7;
		end
		32'h00007550: begin
				q			<=			16'h0793;
		end
		32'h00007552: begin
				q			<=			16'h05B7;
		end
		32'h00007554: begin
				q			<=			16'hF06F;
		end
		32'h00007556: begin
				q			<=			16'hF55F;
		end
		32'h00007558: begin
				q			<=			16'h0793;
		end
		32'h0000755A: begin
				q			<=			16'h0540;
		end
		32'h0000755C: begin
				q			<=			16'hE863;
		end
		32'h0000755E: begin
				q			<=			16'h00E7;
		end
		32'h00007560: begin
				q			<=			16'hD793;
		end
		32'h00007562: begin
				q			<=			16'h00C4;
		end
		32'h00007564: begin
				q			<=			16'h8793;
		end
		32'h00007566: begin
				q			<=			16'h06E7;
		end
		32'h00007568: begin
				q			<=			16'hF06F;
		end
		32'h0000756A: begin
				q			<=			16'hF41F;
		end
		32'h0000756C: begin
				q			<=			16'h0793;
		end
		32'h0000756E: begin
				q			<=			16'h1540;
		end
		32'h00007570: begin
				q			<=			16'hE863;
		end
		32'h00007572: begin
				q			<=			16'h00E7;
		end
		32'h00007574: begin
				q			<=			16'hD793;
		end
		32'h00007576: begin
				q			<=			16'h00F4;
		end
		32'h00007578: begin
				q			<=			16'h8793;
		end
		32'h0000757A: begin
				q			<=			16'h0777;
		end
		32'h0000757C: begin
				q			<=			16'hF06F;
		end
		32'h0000757E: begin
				q			<=			16'hF2DF;
		end
		32'h00007580: begin
				q			<=			16'h0693;
		end
		32'h00007582: begin
				q			<=			16'h5540;
		end
		32'h00007584: begin
				q			<=			16'h0793;
		end
		32'h00007586: begin
				q			<=			16'h07E0;
		end
		32'h00007588: begin
				q			<=			16'hE0E3;
		end
		32'h0000758A: begin
				q			<=			16'hF2E6;
		end
		32'h0000758C: begin
				q			<=			16'hD793;
		end
		32'h0000758E: begin
				q			<=			16'h0124;
		end
		32'h00007590: begin
				q			<=			16'h8793;
		end
		32'h00007592: begin
				q			<=			16'h07C7;
		end
		32'h00007594: begin
				q			<=			16'hF06F;
		end
		32'h00007596: begin
				q			<=			16'hF15F;
		end
		32'h00007598: begin
				q			<=			16'h2683;
		end
		32'h0000759A: begin
				q			<=			16'h00C4;
		end
		32'h0000759C: begin
				q			<=			16'h4C63;
		end
		32'h0000759E: begin
				q			<=			16'h0006;
		end
		32'h000075A0: begin
				q			<=			16'h2783;
		end
		32'h000075A2: begin
				q			<=			16'h0084;
		end
		32'h000075A4: begin
				q			<=			16'hA623;
		end
		32'h000075A6: begin
				q			<=			16'h00D7;
		end
		32'h000075A8: begin
				q			<=			16'hA423;
		end
		32'h000075AA: begin
				q			<=			16'h00F6;
		end
		32'h000075AC: begin
				q			<=			16'h07B3;
		end
		32'h000075AE: begin
				q			<=			16'h00E4;
		end
		32'h000075B0: begin
				q			<=			16'hF06F;
		end
		32'h000075B2: begin
				q			<=			16'hECDF;
		end
		32'h000075B4: begin
				q			<=			16'h8413;
		end
		32'h000075B6: begin
				q			<=			16'h0006;
		end
		32'h000075B8: begin
				q			<=			16'hF06F;
		end
		32'h000075BA: begin
				q			<=			16'hF09F;
		end
		32'h000075BC: begin
				q			<=			16'h9697;
		end
		32'h000075BE: begin
				q			<=			16'h0000;
		end
		32'h000075C0: begin
				q			<=			16'hAC23;
		end
		32'h000075C2: begin
				q			<=			16'hDAB6;
		end
		32'h000075C4: begin
				q			<=			16'h9697;
		end
		32'h000075C6: begin
				q			<=			16'h0000;
		end
		32'h000075C8: begin
				q			<=			16'hA623;
		end
		32'h000075CA: begin
				q			<=			16'hDAB6;
		end
		32'h000075CC: begin
				q			<=			16'h4C63;
		end
		32'h000075CE: begin
				q			<=			16'h0006;
		end
		32'h000075D0: begin
				q			<=			16'h0733;
		end
		32'h000075D2: begin
				q			<=			16'h00E4;
		end
		32'h000075D4: begin
				q			<=			16'h2783;
		end
		32'h000075D6: begin
				q			<=			16'h0047;
		end
		32'h000075D8: begin
				q			<=			16'hE793;
		end
		32'h000075DA: begin
				q			<=			16'h0017;
		end
		32'h000075DC: begin
				q			<=			16'h2223;
		end
		32'h000075DE: begin
				q			<=			16'h00F7;
		end
		32'h000075E0: begin
				q			<=			16'hF06F;
		end
		32'h000075E2: begin
				q			<=			16'hF55F;
		end
		32'h000075E4: begin
				q			<=			16'h0693;
		end
		32'h000075E6: begin
				q			<=			16'h1FF0;
		end
		32'h000075E8: begin
				q			<=			16'hA803;
		end
		32'h000075EA: begin
				q			<=			16'h0049;
		end
		32'h000075EC: begin
				q			<=			16'hE263;
		end
		32'h000075EE: begin
				q			<=			16'h1AE6;
		end
		32'h000075F0: begin
				q			<=			16'h5713;
		end
		32'h000075F2: begin
				q			<=			16'h0037;
		end
		32'h000075F4: begin
				q			<=			16'h5613;
		end
		32'h000075F6: begin
				q			<=			16'h4027;
		end
		32'h000075F8: begin
				q			<=			16'h0693;
		end
		32'h000075FA: begin
				q			<=			16'h0010;
		end
		32'h000075FC: begin
				q			<=			16'h0713;
		end
		32'h000075FE: begin
				q			<=			16'h0017;
		end
		32'h00007600: begin
				q			<=			16'h96B3;
		end
		32'h00007602: begin
				q			<=			16'h00C6;
		end
		32'h00007604: begin
				q			<=			16'h1713;
		end
		32'h00007606: begin
				q			<=			16'h0037;
		end
		32'h00007608: begin
				q			<=			16'h8733;
		end
		32'h0000760A: begin
				q			<=			16'h00E9;
		end
		32'h0000760C: begin
				q			<=			16'hE6B3;
		end
		32'h0000760E: begin
				q			<=			16'h0106;
		end
		32'h00007610: begin
				q			<=			16'h9617;
		end
		32'h00007612: begin
				q			<=			16'h0000;
		end
		32'h00007614: begin
				q			<=			16'h2A23;
		end
		32'h00007616: begin
				q			<=			16'hD4D6;
		end
		32'h00007618: begin
				q			<=			16'h2683;
		end
		32'h0000761A: begin
				q			<=			16'h0007;
		end
		32'h0000761C: begin
				q			<=			16'h0613;
		end
		32'h0000761E: begin
				q			<=			16'hFF87;
		end
		32'h00007620: begin
				q			<=			16'h2623;
		end
		32'h00007622: begin
				q			<=			16'h00C4;
		end
		32'h00007624: begin
				q			<=			16'h2423;
		end
		32'h00007626: begin
				q			<=			16'h00D4;
		end
		32'h00007628: begin
				q			<=			16'h2023;
		end
		32'h0000762A: begin
				q			<=			16'h0087;
		end
		32'h0000762C: begin
				q			<=			16'hA623;
		end
		32'h0000762E: begin
				q			<=			16'h0086;
		end
		32'h00007630: begin
				q			<=			16'hD713;
		end
		32'h00007632: begin
				q			<=			16'h4027;
		end
		32'h00007634: begin
				q			<=			16'h0313;
		end
		32'h00007636: begin
				q			<=			16'h0010;
		end
		32'h00007638: begin
				q			<=			16'h1333;
		end
		32'h0000763A: begin
				q			<=			16'h00E3;
		end
		32'h0000763C: begin
				q			<=			16'hA703;
		end
		32'h0000763E: begin
				q			<=			16'h0049;
		end
		32'h00007640: begin
				q			<=			16'h6C63;
		end
		32'h00007642: begin
				q			<=			16'h0667;
		end
		32'h00007644: begin
				q			<=			16'h76B3;
		end
		32'h00007646: begin
				q			<=			16'h0067;
		end
		32'h00007648: begin
				q			<=			16'h9C63;
		end
		32'h0000764A: begin
				q			<=			16'h0006;
		end
		32'h0000764C: begin
				q			<=			16'hF793;
		end
		32'h0000764E: begin
				q			<=			16'hFFC7;
		end
		32'h00007650: begin
				q			<=			16'h1313;
		end
		32'h00007652: begin
				q			<=			16'h0013;
		end
		32'h00007654: begin
				q			<=			16'h76B3;
		end
		32'h00007656: begin
				q			<=			16'h0067;
		end
		32'h00007658: begin
				q			<=			16'h8793;
		end
		32'h0000765A: begin
				q			<=			16'h0047;
		end
		32'h0000765C: begin
				q			<=			16'h8AE3;
		end
		32'h0000765E: begin
				q			<=			16'hFE06;
		end
		32'h00007660: begin
				q			<=			16'h0E13;
		end
		32'h00007662: begin
				q			<=			16'h00F0;
		end
		32'h00007664: begin
				q			<=			16'h9693;
		end
		32'h00007666: begin
				q			<=			16'h0037;
		end
		32'h00007668: begin
				q			<=			16'h86B3;
		end
		32'h0000766A: begin
				q			<=			16'h00D9;
		end
		32'h0000766C: begin
				q			<=			16'h8813;
		end
		32'h0000766E: begin
				q			<=			16'h0006;
		end
		32'h00007670: begin
				q			<=			16'h8513;
		end
		32'h00007672: begin
				q			<=			16'h0007;
		end
		32'h00007674: begin
				q			<=			16'h2403;
		end
		32'h00007676: begin
				q			<=			16'h00C8;
		end
		32'h00007678: begin
				q			<=			16'h1E63;
		end
		32'h0000767A: begin
				q			<=			16'h1D04;
		end
		32'h0000767C: begin
				q			<=			16'h0513;
		end
		32'h0000767E: begin
				q			<=			16'h0015;
		end
		32'h00007680: begin
				q			<=			16'h7713;
		end
		32'h00007682: begin
				q			<=			16'h0035;
		end
		32'h00007684: begin
				q			<=			16'h0813;
		end
		32'h00007686: begin
				q			<=			16'h0088;
		end
		32'h00007688: begin
				q			<=			16'h16E3;
		end
		32'h0000768A: begin
				q			<=			16'hFE07;
		end
		32'h0000768C: begin
				q			<=			16'hF713;
		end
		32'h0000768E: begin
				q			<=			16'h0037;
		end
		32'h00007690: begin
				q			<=			16'h1463;
		end
		32'h00007692: begin
				q			<=			16'h2407;
		end
		32'h00007694: begin
				q			<=			16'hA703;
		end
		32'h00007696: begin
				q			<=			16'h0049;
		end
		32'h00007698: begin
				q			<=			16'h4793;
		end
		32'h0000769A: begin
				q			<=			16'hFFF3;
		end
		32'h0000769C: begin
				q			<=			16'h77B3;
		end
		32'h0000769E: begin
				q			<=			16'h00F7;
		end
		32'h000076A0: begin
				q			<=			16'h9717;
		end
		32'h000076A2: begin
				q			<=			16'h0000;
		end
		32'h000076A4: begin
				q			<=			16'h2223;
		end
		32'h000076A6: begin
				q			<=			16'hCCF7;
		end
		32'h000076A8: begin
				q			<=			16'hA703;
		end
		32'h000076AA: begin
				q			<=			16'h0049;
		end
		32'h000076AC: begin
				q			<=			16'h1313;
		end
		32'h000076AE: begin
				q			<=			16'h0013;
		end
		32'h000076B0: begin
				q			<=			16'h6463;
		end
		32'h000076B2: begin
				q			<=			16'h0067;
		end
		32'h000076B4: begin
				q			<=			16'h1663;
		end
		32'h000076B6: begin
				q			<=			16'h2403;
		end
		32'h000076B8: begin
				q			<=			16'hAB83;
		end
		32'h000076BA: begin
				q			<=			16'h0089;
		end
		32'h000076BC: begin
				q			<=			16'hA403;
		end
		32'h000076BE: begin
				q			<=			16'h004B;
		end
		32'h000076C0: begin
				q			<=			16'h7A93;
		end
		32'h000076C2: begin
				q			<=			16'hFFC4;
		end
		32'h000076C4: begin
				q			<=			16'hE863;
		end
		32'h000076C6: begin
				q			<=			16'h009A;
		end
		32'h000076C8: begin
				q			<=			16'h8733;
		end
		32'h000076CA: begin
				q			<=			16'h409A;
		end
		32'h000076CC: begin
				q			<=			16'h0793;
		end
		32'h000076CE: begin
				q			<=			16'h00F0;
		end
		32'h000076D0: begin
				q			<=			16'hC463;
		end
		32'h000076D2: begin
				q			<=			16'h36E7;
		end
		32'h000076D4: begin
				q			<=			16'hA797;
		end
		32'h000076D6: begin
				q			<=			16'h0000;
		end
		32'h000076D8: begin
				q			<=			16'h8793;
		end
		32'h000076DA: begin
				q			<=			16'h8D47;
		end
		32'h000076DC: begin
				q			<=			16'hA403;
		end
		32'h000076DE: begin
				q			<=			16'h0007;
		end
		32'h000076E0: begin
				q			<=			16'h9797;
		end
		32'h000076E2: begin
				q			<=			16'h0000;
		end
		32'h000076E4: begin
				q			<=			16'h8793;
		end
		32'h000076E6: begin
				q			<=			16'h1FC7;
		end
		32'h000076E8: begin
				q			<=			16'hA683;
		end
		32'h000076EA: begin
				q			<=			16'h0007;
		end
		32'h000076EC: begin
				q			<=			16'h0713;
		end
		32'h000076EE: begin
				q			<=			16'hFFF0;
		end
		32'h000076F0: begin
				q			<=			16'h8433;
		end
		32'h000076F2: begin
				q			<=			16'h0084;
		end
		32'h000076F4: begin
				q			<=			16'h8A13;
		end
		32'h000076F6: begin
				q			<=			16'h0007;
		end
		32'h000076F8: begin
				q			<=			16'h9863;
		end
		32'h000076FA: begin
				q			<=			16'h20E6;
		end
		32'h000076FC: begin
				q			<=			16'h0413;
		end
		32'h000076FE: begin
				q			<=			16'h0104;
		end
		32'h00007700: begin
				q			<=			16'h0593;
		end
		32'h00007702: begin
				q			<=			16'h0004;
		end
		32'h00007704: begin
				q			<=			16'h0513;
		end
		32'h00007706: begin
				q			<=			16'h0009;
		end
		32'h00007708: begin
				q			<=			16'h10EF;
		end
		32'h0000770A: begin
				q			<=			16'h3000;
		end
		32'h0000770C: begin
				q			<=			16'h0793;
		end
		32'h0000770E: begin
				q			<=			16'hFFF0;
		end
		32'h00007710: begin
				q			<=			16'h0B13;
		end
		32'h00007712: begin
				q			<=			16'h0005;
		end
		32'h00007714: begin
				q			<=			16'h0263;
		end
		32'h00007716: begin
				q			<=			16'h2AF5;
		end
		32'h00007718: begin
				q			<=			16'h87B3;
		end
		32'h0000771A: begin
				q			<=			16'h015B;
		end
		32'h0000771C: begin
				q			<=			16'h7463;
		end
		32'h0000771E: begin
				q			<=			16'h00F5;
		end
		32'h00007720: begin
				q			<=			16'h9C63;
		end
		32'h00007722: begin
				q			<=			16'h293B;
		end
		32'h00007724: begin
				q			<=			16'h9C17;
		end
		32'h00007726: begin
				q			<=			16'h0000;
		end
		32'h00007728: begin
				q			<=			16'h0C13;
		end
		32'h0000772A: begin
				q			<=			16'h3D0C;
		end
		32'h0000772C: begin
				q			<=			16'h2703;
		end
		32'h0000772E: begin
				q			<=			16'h000C;
		end
		32'h00007730: begin
				q			<=			16'h0733;
		end
		32'h00007732: begin
				q			<=			16'h00E4;
		end
		32'h00007734: begin
				q			<=			16'h9697;
		end
		32'h00007736: begin
				q			<=			16'h0000;
		end
		32'h00007738: begin
				q			<=			16'hA023;
		end
		32'h0000773A: begin
				q			<=			16'h3CE6;
		end
		32'h0000773C: begin
				q			<=			16'h9263;
		end
		32'h0000773E: begin
				q			<=			16'h1F67;
		end
		32'h00007740: begin
				q			<=			16'h9693;
		end
		32'h00007742: begin
				q			<=			16'h0147;
		end
		32'h00007744: begin
				q			<=			16'h9E63;
		end
		32'h00007746: begin
				q			<=			16'h1C06;
		end
		32'h00007748: begin
				q			<=			16'hA783;
		end
		32'h0000774A: begin
				q			<=			16'h0089;
		end
		32'h0000774C: begin
				q			<=			16'h8433;
		end
		32'h0000774E: begin
				q			<=			16'h008A;
		end
		32'h00007750: begin
				q			<=			16'h6413;
		end
		32'h00007752: begin
				q			<=			16'h0014;
		end
		32'h00007754: begin
				q			<=			16'hA223;
		end
		32'h00007756: begin
				q			<=			16'h0087;
		end
		32'h00007758: begin
				q			<=			16'hA717;
		end
		32'h0000775A: begin
				q			<=			16'h0000;
		end
		32'h0000775C: begin
				q			<=			16'h0713;
		end
		32'h0000775E: begin
				q			<=			16'h84C7;
		end
		32'h00007760: begin
				q			<=			16'h2783;
		end
		32'h00007762: begin
				q			<=			16'h000C;
		end
		32'h00007764: begin
				q			<=			16'h2703;
		end
		32'h00007766: begin
				q			<=			16'h0007;
		end
		32'h00007768: begin
				q			<=			16'h7663;
		end
		32'h0000776A: begin
				q			<=			16'h00F7;
		end
		32'h0000776C: begin
				q			<=			16'hA717;
		end
		32'h0000776E: begin
				q			<=			16'h0000;
		end
		32'h00007770: begin
				q			<=			16'h2C23;
		end
		32'h00007772: begin
				q			<=			16'h82F7;
		end
		32'h00007774: begin
				q			<=			16'hA717;
		end
		32'h00007776: begin
				q			<=			16'h0000;
		end
		32'h00007778: begin
				q			<=			16'h0713;
		end
		32'h0000777A: begin
				q			<=			16'h82C7;
		end
		32'h0000777C: begin
				q			<=			16'h2703;
		end
		32'h0000777E: begin
				q			<=			16'h0007;
		end
		32'h00007780: begin
				q			<=			16'h7C63;
		end
		32'h00007782: begin
				q			<=			16'h22F7;
		end
		32'h00007784: begin
				q			<=			16'hA717;
		end
		32'h00007786: begin
				q			<=			16'h0000;
		end
		32'h00007788: begin
				q			<=			16'h2E23;
		end
		32'h0000778A: begin
				q			<=			16'h80F7;
		end
		32'h0000778C: begin
				q			<=			16'h006F;
		end
		32'h0000778E: begin
				q			<=			16'h22C0;
		end
		32'h00007790: begin
				q			<=			16'h5613;
		end
		32'h00007792: begin
				q			<=			16'h0097;
		end
		32'h00007794: begin
				q			<=			16'h0693;
		end
		32'h00007796: begin
				q			<=			16'h0040;
		end
		32'h00007798: begin
				q			<=			16'hE863;
		end
		32'h0000779A: begin
				q			<=			16'h04C6;
		end
		32'h0000779C: begin
				q			<=			16'h5693;
		end
		32'h0000779E: begin
				q			<=			16'h0067;
		end
		32'h000077A0: begin
				q			<=			16'h8693;
		end
		32'h000077A2: begin
				q			<=			16'h0386;
		end
		32'h000077A4: begin
				q			<=			16'h8613;
		end
		32'h000077A6: begin
				q			<=			16'h0016;
		end
		32'h000077A8: begin
				q			<=			16'h1613;
		end
		32'h000077AA: begin
				q			<=			16'h0036;
		end
		32'h000077AC: begin
				q			<=			16'h8633;
		end
		32'h000077AE: begin
				q			<=			16'h00C9;
		end
		32'h000077B0: begin
				q			<=			16'h0513;
		end
		32'h000077B2: begin
				q			<=			16'hFF86;
		end
		32'h000077B4: begin
				q			<=			16'h2603;
		end
		32'h000077B6: begin
				q			<=			16'h0006;
		end
		32'h000077B8: begin
				q			<=			16'h1463;
		end
		32'h000077BA: begin
				q			<=			16'h08C5;
		end
		32'h000077BC: begin
				q			<=			16'h0713;
		end
		32'h000077BE: begin
				q			<=			16'h0010;
		end
		32'h000077C0: begin
				q			<=			16'hD693;
		end
		32'h000077C2: begin
				q			<=			16'h4026;
		end
		32'h000077C4: begin
				q			<=			16'h16B3;
		end
		32'h000077C6: begin
				q			<=			16'h00D7;
		end
		32'h000077C8: begin
				q			<=			16'hE6B3;
		end
		32'h000077CA: begin
				q			<=			16'h0106;
		end
		32'h000077CC: begin
				q			<=			16'h9717;
		end
		32'h000077CE: begin
				q			<=			16'h0000;
		end
		32'h000077D0: begin
				q			<=			16'h2C23;
		end
		32'h000077D2: begin
				q			<=			16'hB8D7;
		end
		32'h000077D4: begin
				q			<=			16'h2623;
		end
		32'h000077D6: begin
				q			<=			16'h00A4;
		end
		32'h000077D8: begin
				q			<=			16'h2423;
		end
		32'h000077DA: begin
				q			<=			16'h00C4;
		end
		32'h000077DC: begin
				q			<=			16'h2423;
		end
		32'h000077DE: begin
				q			<=			16'h0085;
		end
		32'h000077E0: begin
				q			<=			16'h2623;
		end
		32'h000077E2: begin
				q			<=			16'h0086;
		end
		32'h000077E4: begin
				q			<=			16'hF06F;
		end
		32'h000077E6: begin
				q			<=			16'hE4DF;
		end
		32'h000077E8: begin
				q			<=			16'h0693;
		end
		32'h000077EA: begin
				q			<=			16'h0140;
		end
		32'h000077EC: begin
				q			<=			16'hE663;
		end
		32'h000077EE: begin
				q			<=			16'h00C6;
		end
		32'h000077F0: begin
				q			<=			16'h0693;
		end
		32'h000077F2: begin
				q			<=			16'h05B6;
		end
		32'h000077F4: begin
				q			<=			16'hF06F;
		end
		32'h000077F6: begin
				q			<=			16'hFB1F;
		end
		32'h000077F8: begin
				q			<=			16'h0693;
		end
		32'h000077FA: begin
				q			<=			16'h0540;
		end
		32'h000077FC: begin
				q			<=			16'hE863;
		end
		32'h000077FE: begin
				q			<=			16'h00C6;
		end
		32'h00007800: begin
				q			<=			16'h5693;
		end
		32'h00007802: begin
				q			<=			16'h00C7;
		end
		32'h00007804: begin
				q			<=			16'h8693;
		end
		32'h00007806: begin
				q			<=			16'h06E6;
		end
		32'h00007808: begin
				q			<=			16'hF06F;
		end
		32'h0000780A: begin
				q			<=			16'hF9DF;
		end
		32'h0000780C: begin
				q			<=			16'h0693;
		end
		32'h0000780E: begin
				q			<=			16'h1540;
		end
		32'h00007810: begin
				q			<=			16'hE863;
		end
		32'h00007812: begin
				q			<=			16'h00C6;
		end
		32'h00007814: begin
				q			<=			16'h5693;
		end
		32'h00007816: begin
				q			<=			16'h00F7;
		end
		32'h00007818: begin
				q			<=			16'h8693;
		end
		32'h0000781A: begin
				q			<=			16'h0776;
		end
		32'h0000781C: begin
				q			<=			16'hF06F;
		end
		32'h0000781E: begin
				q			<=			16'hF89F;
		end
		32'h00007820: begin
				q			<=			16'h0513;
		end
		32'h00007822: begin
				q			<=			16'h5540;
		end
		32'h00007824: begin
				q			<=			16'h0693;
		end
		32'h00007826: begin
				q			<=			16'h07E0;
		end
		32'h00007828: begin
				q			<=			16'h6EE3;
		end
		32'h0000782A: begin
				q			<=			16'hF6C5;
		end
		32'h0000782C: begin
				q			<=			16'h5693;
		end
		32'h0000782E: begin
				q			<=			16'h0127;
		end
		32'h00007830: begin
				q			<=			16'h8693;
		end
		32'h00007832: begin
				q			<=			16'h07C6;
		end
		32'h00007834: begin
				q			<=			16'hF06F;
		end
		32'h00007836: begin
				q			<=			16'hF71F;
		end
		32'h00007838: begin
				q			<=			16'h2603;
		end
		32'h0000783A: begin
				q			<=			16'h0086;
		end
		32'h0000783C: begin
				q			<=			16'h0863;
		end
		32'h0000783E: begin
				q			<=			16'h00C5;
		end
		32'h00007840: begin
				q			<=			16'h2683;
		end
		32'h00007842: begin
				q			<=			16'h0046;
		end
		32'h00007844: begin
				q			<=			16'hF693;
		end
		32'h00007846: begin
				q			<=			16'hFFC6;
		end
		32'h00007848: begin
				q			<=			16'h68E3;
		end
		32'h0000784A: begin
				q			<=			16'hFED7;
		end
		32'h0000784C: begin
				q			<=			16'h2503;
		end
		32'h0000784E: begin
				q			<=			16'h00C6;
		end
		32'h00007850: begin
				q			<=			16'hF06F;
		end
		32'h00007852: begin
				q			<=			16'hF85F;
		end
		32'h00007854: begin
				q			<=			16'h2703;
		end
		32'h00007856: begin
				q			<=			16'h0044;
		end
		32'h00007858: begin
				q			<=			16'h2603;
		end
		32'h0000785A: begin
				q			<=			16'h00C4;
		end
		32'h0000785C: begin
				q			<=			16'h7713;
		end
		32'h0000785E: begin
				q			<=			16'hFFC7;
		end
		32'h00007860: begin
				q			<=			16'h08B3;
		end
		32'h00007862: begin
				q			<=			16'h4097;
		end
		32'h00007864: begin
				q			<=			16'h5463;
		end
		32'h00007866: begin
				q			<=			16'h051E;
		end
		32'h00007868: begin
				q			<=			16'hE793;
		end
		32'h0000786A: begin
				q			<=			16'h0014;
		end
		32'h0000786C: begin
				q			<=			16'h2223;
		end
		32'h0000786E: begin
				q			<=			16'h00F4;
		end
		32'h00007870: begin
				q			<=			16'h2783;
		end
		32'h00007872: begin
				q			<=			16'h0084;
		end
		32'h00007874: begin
				q			<=			16'h06B3;
		end
		32'h00007876: begin
				q			<=			16'h0094;
		end
		32'h00007878: begin
				q			<=			16'h0733;
		end
		32'h0000787A: begin
				q			<=			16'h00E4;
		end
		32'h0000787C: begin
				q			<=			16'hA623;
		end
		32'h0000787E: begin
				q			<=			16'h00C7;
		end
		32'h00007880: begin
				q			<=			16'h2423;
		end
		32'h00007882: begin
				q			<=			16'h00F6;
		end
		32'h00007884: begin
				q			<=			16'h9797;
		end
		32'h00007886: begin
				q			<=			16'h0000;
		end
		32'h00007888: begin
				q			<=			16'hA823;
		end
		32'h0000788A: begin
				q			<=			16'hAED7;
		end
		32'h0000788C: begin
				q			<=			16'h9797;
		end
		32'h0000788E: begin
				q			<=			16'h0000;
		end
		32'h00007890: begin
				q			<=			16'hA223;
		end
		32'h00007892: begin
				q			<=			16'hAED7;
		end
		32'h00007894: begin
				q			<=			16'hE793;
		end
		32'h00007896: begin
				q			<=			16'h0018;
		end
		32'h00007898: begin
				q			<=			16'hA623;
		end
		32'h0000789A: begin
				q			<=			16'h00B6;
		end
		32'h0000789C: begin
				q			<=			16'hA423;
		end
		32'h0000789E: begin
				q			<=			16'h00B6;
		end
		32'h000078A0: begin
				q			<=			16'hA223;
		end
		32'h000078A2: begin
				q			<=			16'h00F6;
		end
		32'h000078A4: begin
				q			<=			16'h2023;
		end
		32'h000078A6: begin
				q			<=			16'h0117;
		end
		32'h000078A8: begin
				q			<=			16'hF06F;
		end
		32'h000078AA: begin
				q			<=			16'hC8DF;
		end
		32'h000078AC: begin
				q			<=			16'hC263;
		end
		32'h000078AE: begin
				q			<=			16'h0208;
		end
		32'h000078B0: begin
				q			<=			16'h0733;
		end
		32'h000078B2: begin
				q			<=			16'h00E4;
		end
		32'h000078B4: begin
				q			<=			16'h2783;
		end
		32'h000078B6: begin
				q			<=			16'h0047;
		end
		32'h000078B8: begin
				q			<=			16'hE793;
		end
		32'h000078BA: begin
				q			<=			16'h0017;
		end
		32'h000078BC: begin
				q			<=			16'h2223;
		end
		32'h000078BE: begin
				q			<=			16'h00F7;
		end
		32'h000078C0: begin
				q			<=			16'h2783;
		end
		32'h000078C2: begin
				q			<=			16'h0084;
		end
		32'h000078C4: begin
				q			<=			16'hA623;
		end
		32'h000078C6: begin
				q			<=			16'h00C7;
		end
		32'h000078C8: begin
				q			<=			16'h2423;
		end
		32'h000078CA: begin
				q			<=			16'h00F6;
		end
		32'h000078CC: begin
				q			<=			16'hF06F;
		end
		32'h000078CE: begin
				q			<=			16'hC69F;
		end
		32'h000078D0: begin
				q			<=			16'h0413;
		end
		32'h000078D2: begin
				q			<=			16'h0006;
		end
		32'h000078D4: begin
				q			<=			16'hF06F;
		end
		32'h000078D6: begin
				q			<=			16'hDA5F;
		end
		32'h000078D8: begin
				q			<=			16'h8713;
		end
		32'h000078DA: begin
				q			<=			16'hFF86;
		end
		32'h000078DC: begin
				q			<=			16'hA683;
		end
		32'h000078DE: begin
				q			<=			16'h0006;
		end
		32'h000078E0: begin
				q			<=			16'h8793;
		end
		32'h000078E2: begin
				q			<=			16'hFFF7;
		end
		32'h000078E4: begin
				q			<=			16'h84E3;
		end
		32'h000078E6: begin
				q			<=			16'hDAE6;
		end
		32'h000078E8: begin
				q			<=			16'hF06F;
		end
		32'h000078EA: begin
				q			<=			16'hDC1F;
		end
		32'h000078EC: begin
				q			<=			16'h8793;
		end
		32'h000078EE: begin
				q			<=			16'h0047;
		end
		32'h000078F0: begin
				q			<=			16'h1313;
		end
		32'h000078F2: begin
				q			<=			16'h0013;
		end
		32'h000078F4: begin
				q			<=			16'h76B3;
		end
		32'h000078F6: begin
				q			<=			16'h0067;
		end
		32'h000078F8: begin
				q			<=			16'h8AE3;
		end
		32'h000078FA: begin
				q			<=			16'hFE06;
		end
		32'h000078FC: begin
				q			<=			16'hF06F;
		end
		32'h000078FE: begin
				q			<=			16'hD69F;
		end
		32'h00007900: begin
				q			<=			16'h0793;
		end
		32'h00007902: begin
				q			<=			16'h0005;
		end
		32'h00007904: begin
				q			<=			16'hF06F;
		end
		32'h00007906: begin
				q			<=			16'hFF1F;
		end
		32'h00007908: begin
				q			<=			16'h17B7;
		end
		32'h0000790A: begin
				q			<=			16'h0000;
		end
		32'h0000790C: begin
				q			<=			16'h8793;
		end
		32'h0000790E: begin
				q			<=			16'h00F7;
		end
		32'h00007910: begin
				q			<=			16'h0433;
		end
		32'h00007912: begin
				q			<=			16'h00F4;
		end
		32'h00007914: begin
				q			<=			16'hF7B7;
		end
		32'h00007916: begin
				q			<=			16'hFFFF;
		end
		32'h00007918: begin
				q			<=			16'h7433;
		end
		32'h0000791A: begin
				q			<=			16'h00F4;
		end
		32'h0000791C: begin
				q			<=			16'hF06F;
		end
		32'h0000791E: begin
				q			<=			16'hDE5F;
		end
		32'h00007920: begin
				q			<=			16'h2603;
		end
		32'h00007922: begin
				q			<=			16'h000A;
		end
		32'h00007924: begin
				q			<=			16'h0693;
		end
		32'h00007926: begin
				q			<=			16'hFFF0;
		end
		32'h00007928: begin
				q			<=			16'h1E63;
		end
		32'h0000792A: begin
				q			<=			16'h0AD6;
		end
		32'h0000792C: begin
				q			<=			16'h9797;
		end
		32'h0000792E: begin
				q			<=			16'h0000;
		end
		32'h00007930: begin
				q			<=			16'hA823;
		end
		32'h00007932: begin
				q			<=			16'hFB67;
		end
		32'h00007934: begin
				q			<=			16'h7593;
		end
		32'h00007936: begin
				q			<=			16'h007B;
		end
		32'h00007938: begin
				q			<=			16'h8863;
		end
		32'h0000793A: begin
				q			<=			16'h0005;
		end
		32'h0000793C: begin
				q			<=			16'h0793;
		end
		32'h0000793E: begin
				q			<=			16'h0080;
		end
		32'h00007940: begin
				q			<=			16'h85B3;
		end
		32'h00007942: begin
				q			<=			16'h40B7;
		end
		32'h00007944: begin
				q			<=			16'h0B33;
		end
		32'h00007946: begin
				q			<=			16'h00BB;
		end
		32'h00007948: begin
				q			<=			16'h17B7;
		end
		32'h0000794A: begin
				q			<=			16'h0000;
		end
		32'h0000794C: begin
				q			<=			16'h85B3;
		end
		32'h0000794E: begin
				q			<=			16'h00F5;
		end
		32'h00007950: begin
				q			<=			16'h0433;
		end
		32'h00007952: begin
				q			<=			16'h008B;
		end
		32'h00007954: begin
				q			<=			16'h8793;
		end
		32'h00007956: begin
				q			<=			16'hFFF7;
		end
		32'h00007958: begin
				q			<=			16'h7433;
		end
		32'h0000795A: begin
				q			<=			16'h00F4;
		end
		32'h0000795C: begin
				q			<=			16'h8A33;
		end
		32'h0000795E: begin
				q			<=			16'h4085;
		end
		32'h00007960: begin
				q			<=			16'h0593;
		end
		32'h00007962: begin
				q			<=			16'h000A;
		end
		32'h00007964: begin
				q			<=			16'h0513;
		end
		32'h00007966: begin
				q			<=			16'h0009;
		end
		32'h00007968: begin
				q			<=			16'h10EF;
		end
		32'h0000796A: begin
				q			<=			16'h0A00;
		end
		32'h0000796C: begin
				q			<=			16'h0793;
		end
		32'h0000796E: begin
				q			<=			16'hFFF0;
		end
		32'h00007970: begin
				q			<=			16'h1663;
		end
		32'h00007972: begin
				q			<=			16'h00F5;
		end
		32'h00007974: begin
				q			<=			16'h0513;
		end
		32'h00007976: begin
				q			<=			16'h000B;
		end
		32'h00007978: begin
				q			<=			16'h0A13;
		end
		32'h0000797A: begin
				q			<=			16'h0000;
		end
		32'h0000797C: begin
				q			<=			16'h2783;
		end
		32'h0000797E: begin
				q			<=			16'h000C;
		end
		32'h00007980: begin
				q			<=			16'h0533;
		end
		32'h00007982: begin
				q			<=			16'h4165;
		end
		32'h00007984: begin
				q			<=			16'h87B3;
		end
		32'h00007986: begin
				q			<=			16'h0147;
		end
		32'h00007988: begin
				q			<=			16'h0A33;
		end
		32'h0000798A: begin
				q			<=			16'h0145;
		end
		32'h0000798C: begin
				q			<=			16'h9717;
		end
		32'h0000798E: begin
				q			<=			16'h0000;
		end
		32'h00007990: begin
				q			<=			16'h2423;
		end
		32'h00007992: begin
				q			<=			16'h16F7;
		end
		32'h00007994: begin
				q			<=			16'h6A13;
		end
		32'h00007996: begin
				q			<=			16'h001A;
		end
		32'h00007998: begin
				q			<=			16'h9797;
		end
		32'h0000799A: begin
				q			<=			16'h0000;
		end
		32'h0000799C: begin
				q			<=			16'hA823;
		end
		32'h0000799E: begin
				q			<=			16'h9D67;
		end
		32'h000079A0: begin
				q			<=			16'h2223;
		end
		32'h000079A2: begin
				q			<=			16'h014B;
		end
		32'h000079A4: begin
				q			<=			16'h8AE3;
		end
		32'h000079A6: begin
				q			<=			16'hDB3B;
		end
		32'h000079A8: begin
				q			<=			16'h0713;
		end
		32'h000079AA: begin
				q			<=			16'h00F0;
		end
		32'h000079AC: begin
				q			<=			16'h6663;
		end
		32'h000079AE: begin
				q			<=			16'h0557;
		end
		32'h000079B0: begin
				q			<=			16'h0793;
		end
		32'h000079B2: begin
				q			<=			16'h0010;
		end
		32'h000079B4: begin
				q			<=			16'h2223;
		end
		32'h000079B6: begin
				q			<=			16'h00FB;
		end
		32'h000079B8: begin
				q			<=			16'hA783;
		end
		32'h000079BA: begin
				q			<=			16'h0089;
		end
		32'h000079BC: begin
				q			<=			16'hA783;
		end
		32'h000079BE: begin
				q			<=			16'h0047;
		end
		32'h000079C0: begin
				q			<=			16'hF793;
		end
		32'h000079C2: begin
				q			<=			16'hFFC7;
		end
		32'h000079C4: begin
				q			<=			16'h8733;
		end
		32'h000079C6: begin
				q			<=			16'h4097;
		end
		32'h000079C8: begin
				q			<=			16'hE663;
		end
		32'h000079CA: begin
				q			<=			16'h0097;
		end
		32'h000079CC: begin
				q			<=			16'h0793;
		end
		32'h000079CE: begin
				q			<=			16'h00F0;
		end
		32'h000079D0: begin
				q			<=			16'hC463;
		end
		32'h000079D2: begin
				q			<=			16'h06E7;
		end
		32'h000079D4: begin
				q			<=			16'h0513;
		end
		32'h000079D6: begin
				q			<=			16'h0009;
		end
		32'h000079D8: begin
				q			<=			16'h0097;
		end
		32'h000079DA: begin
				q			<=			16'h0000;
		end
		32'h000079DC: begin
				q			<=			16'h80E7;
		end
		32'h000079DE: begin
				q			<=			16'h0AC0;
		end
		32'h000079E0: begin
				q			<=			16'hF06F;
		end
		32'h000079E2: begin
				q			<=			16'hA09F;
		end
		32'h000079E4: begin
				q			<=			16'h07B3;
		end
		32'h000079E6: begin
				q			<=			16'h40FB;
		end
		32'h000079E8: begin
				q			<=			16'h87B3;
		end
		32'h000079EA: begin
				q			<=			16'h00E7;
		end
		32'h000079EC: begin
				q			<=			16'h9717;
		end
		32'h000079EE: begin
				q			<=			16'h0000;
		end
		32'h000079F0: begin
				q			<=			16'h2423;
		end
		32'h000079F2: begin
				q			<=			16'h10F7;
		end
		32'h000079F4: begin
				q			<=			16'hF06F;
		end
		32'h000079F6: begin
				q			<=			16'hF41F;
		end
		32'h000079F8: begin
				q			<=			16'hA783;
		end
		32'h000079FA: begin
				q			<=			16'h004B;
		end
		32'h000079FC: begin
				q			<=			16'h8413;
		end
		32'h000079FE: begin
				q			<=			16'hFF4A;
		end
		32'h00007A00: begin
				q			<=			16'h7413;
		end
		32'h00007A02: begin
				q			<=			16'hFF84;
		end
		32'h00007A04: begin
				q			<=			16'hF793;
		end
		32'h00007A06: begin
				q			<=			16'h0017;
		end
		32'h00007A08: begin
				q			<=			16'hE7B3;
		end
		32'h00007A0A: begin
				q			<=			16'h0087;
		end
		32'h00007A0C: begin
				q			<=			16'hA223;
		end
		32'h00007A0E: begin
				q			<=			16'h00FB;
		end
		32'h00007A10: begin
				q			<=			16'h0693;
		end
		32'h00007A12: begin
				q			<=			16'h0050;
		end
		32'h00007A14: begin
				q			<=			16'h87B3;
		end
		32'h00007A16: begin
				q			<=			16'h008B;
		end
		32'h00007A18: begin
				q			<=			16'hA223;
		end
		32'h00007A1A: begin
				q			<=			16'h00D7;
		end
		32'h00007A1C: begin
				q			<=			16'hA423;
		end
		32'h00007A1E: begin
				q			<=			16'h00D7;
		end
		32'h00007A20: begin
				q			<=			16'h7CE3;
		end
		32'h00007A22: begin
				q			<=			16'hD287;
		end
		32'h00007A24: begin
				q			<=			16'h8593;
		end
		32'h00007A26: begin
				q			<=			16'h008B;
		end
		32'h00007A28: begin
				q			<=			16'h0513;
		end
		32'h00007A2A: begin
				q			<=			16'h0009;
		end
		32'h00007A2C: begin
				q			<=			16'hD097;
		end
		32'h00007A2E: begin
				q			<=			16'hFFFF;
		end
		32'h00007A30: begin
				q			<=			16'h80E7;
		end
		32'h00007A32: begin
				q			<=			16'h5440;
		end
		32'h00007A34: begin
				q			<=			16'hF06F;
		end
		32'h00007A36: begin
				q			<=			16'hD25F;
		end
		32'h00007A38: begin
				q			<=			16'hA403;
		end
		32'h00007A3A: begin
				q			<=			16'h0089;
		end
		32'h00007A3C: begin
				q			<=			16'hE793;
		end
		32'h00007A3E: begin
				q			<=			16'h0014;
		end
		32'h00007A40: begin
				q			<=			16'h2223;
		end
		32'h00007A42: begin
				q			<=			16'h00F4;
		end
		32'h00007A44: begin
				q			<=			16'h07B3;
		end
		32'h00007A46: begin
				q			<=			16'h0094;
		end
		32'h00007A48: begin
				q			<=			16'h9697;
		end
		32'h00007A4A: begin
				q			<=			16'h0000;
		end
		32'h00007A4C: begin
				q			<=			16'hA023;
		end
		32'h00007A4E: begin
				q			<=			16'h92F6;
		end
		32'h00007A50: begin
				q			<=			16'hF06F;
		end
		32'h00007A52: begin
				q			<=			16'hA31F;
		end
		32'h00007A54: begin
				q			<=			16'h0000;
		end
		32'h00007A56: begin
				q			<=			16'h0000;
		end
		32'h00007A58: begin
				q			<=			16'hF593;
		end
		32'h00007A5A: begin
				q			<=			16'h0FF5;
		end
		32'h00007A5C: begin
				q			<=			16'h0633;
		end
		32'h00007A5E: begin
				q			<=			16'h00C5;
		end
		32'h00007A60: begin
				q			<=			16'h1663;
		end
		32'h00007A62: begin
				q			<=			16'h00C5;
		end
		32'h00007A64: begin
				q			<=			16'h0513;
		end
		32'h00007A66: begin
				q			<=			16'h0000;
		end
		32'h00007A68: begin
				q			<=			16'h8067;
		end
		32'h00007A6A: begin
				q			<=			16'h0000;
		end
		32'h00007A6C: begin
				q			<=			16'h4783;
		end
		32'h00007A6E: begin
				q			<=			16'h0005;
		end
		32'h00007A70: begin
				q			<=			16'h8CE3;
		end
		32'h00007A72: begin
				q			<=			16'hFEB7;
		end
		32'h00007A74: begin
				q			<=			16'h0513;
		end
		32'h00007A76: begin
				q			<=			16'h0015;
		end
		32'h00007A78: begin
				q			<=			16'hF06F;
		end
		32'h00007A7A: begin
				q			<=			16'hFE9F;
		end
		32'h00007A7C: begin
				q			<=			16'h0000;
		end
		32'h00007A7E: begin
				q			<=			16'h0000;
		end
		32'h00007A80: begin
				q			<=			16'h8067;
		end
		32'h00007A82: begin
				q			<=			16'h0000;
		end
		32'h00007A84: begin
				q			<=			16'h8067;
		end
		32'h00007A86: begin
				q			<=			16'h0000;
		end
		32'h00007A88: begin
				q			<=			16'h0000;
		end
		32'h00007A8A: begin
				q			<=			16'h0000;
		end
		32'h00007A8C: begin
				q			<=			16'h2783;
		end
		32'h00007A8E: begin
				q			<=			16'h04C5;
		end
		32'h00007A90: begin
				q			<=			16'h0113;
		end
		32'h00007A92: begin
				q			<=			16'hFF01;
		end
		32'h00007A94: begin
				q			<=			16'h2223;
		end
		32'h00007A96: begin
				q			<=			16'h0091;
		end
		32'h00007A98: begin
				q			<=			16'h2023;
		end
		32'h00007A9A: begin
				q			<=			16'h0121;
		end
		32'h00007A9C: begin
				q			<=			16'h2623;
		end
		32'h00007A9E: begin
				q			<=			16'h0011;
		end
		32'h00007AA0: begin
				q			<=			16'h2423;
		end
		32'h00007AA2: begin
				q			<=			16'h0081;
		end
		32'h00007AA4: begin
				q			<=			16'h0493;
		end
		32'h00007AA6: begin
				q			<=			16'h0005;
		end
		32'h00007AA8: begin
				q			<=			16'h8913;
		end
		32'h00007AAA: begin
				q			<=			16'h0005;
		end
		32'h00007AAC: begin
				q			<=			16'h8263;
		end
		32'h00007AAE: begin
				q			<=			16'h0407;
		end
		32'h00007AB0: begin
				q			<=			16'hA703;
		end
		32'h00007AB2: begin
				q			<=			16'h04C4;
		end
		32'h00007AB4: begin
				q			<=			16'h1793;
		end
		32'h00007AB6: begin
				q			<=			16'h0029;
		end
		32'h00007AB8: begin
				q			<=			16'h07B3;
		end
		32'h00007ABA: begin
				q			<=			16'h00F7;
		end
		32'h00007ABC: begin
				q			<=			16'hA503;
		end
		32'h00007ABE: begin
				q			<=			16'h0007;
		end
		32'h00007AC0: begin
				q			<=			16'h1063;
		end
		32'h00007AC2: begin
				q			<=			16'h0605;
		end
		32'h00007AC4: begin
				q			<=			16'h0413;
		end
		32'h00007AC6: begin
				q			<=			16'h0010;
		end
		32'h00007AC8: begin
				q			<=			16'h1433;
		end
		32'h00007ACA: begin
				q			<=			16'h0124;
		end
		32'h00007ACC: begin
				q			<=			16'h0613;
		end
		32'h00007ACE: begin
				q			<=			16'h0054;
		end
		32'h00007AD0: begin
				q			<=			16'h1613;
		end
		32'h00007AD2: begin
				q			<=			16'h0026;
		end
		32'h00007AD4: begin
				q			<=			16'h0593;
		end
		32'h00007AD6: begin
				q			<=			16'h0010;
		end
		32'h00007AD8: begin
				q			<=			16'h8513;
		end
		32'h00007ADA: begin
				q			<=			16'h0004;
		end
		32'h00007ADC: begin
				q			<=			16'h10EF;
		end
		32'h00007ADE: begin
				q			<=			16'h6E10;
		end
		32'h00007AE0: begin
				q			<=			16'h0263;
		end
		32'h00007AE2: begin
				q			<=			16'h0205;
		end
		32'h00007AE4: begin
				q			<=			16'h2223;
		end
		32'h00007AE6: begin
				q			<=			16'h0125;
		end
		32'h00007AE8: begin
				q			<=			16'h2423;
		end
		32'h00007AEA: begin
				q			<=			16'h0085;
		end
		32'h00007AEC: begin
				q			<=			16'h006F;
		end
		32'h00007AEE: begin
				q			<=			16'h03C0;
		end
		32'h00007AF0: begin
				q			<=			16'h0613;
		end
		32'h00007AF2: begin
				q			<=			16'h0210;
		end
		32'h00007AF4: begin
				q			<=			16'h0593;
		end
		32'h00007AF6: begin
				q			<=			16'h0040;
		end
		32'h00007AF8: begin
				q			<=			16'h10EF;
		end
		32'h00007AFA: begin
				q			<=			16'h6C50;
		end
		32'h00007AFC: begin
				q			<=			16'hA623;
		end
		32'h00007AFE: begin
				q			<=			16'h04A4;
		end
		32'h00007B00: begin
				q			<=			16'h18E3;
		end
		32'h00007B02: begin
				q			<=			16'hFA05;
		end
		32'h00007B04: begin
				q			<=			16'h0513;
		end
		32'h00007B06: begin
				q			<=			16'h0000;
		end
		32'h00007B08: begin
				q			<=			16'h2083;
		end
		32'h00007B0A: begin
				q			<=			16'h00C1;
		end
		32'h00007B0C: begin
				q			<=			16'h2403;
		end
		32'h00007B0E: begin
				q			<=			16'h0081;
		end
		32'h00007B10: begin
				q			<=			16'h2483;
		end
		32'h00007B12: begin
				q			<=			16'h0041;
		end
		32'h00007B14: begin
				q			<=			16'h2903;
		end
		32'h00007B16: begin
				q			<=			16'h0001;
		end
		32'h00007B18: begin
				q			<=			16'h0113;
		end
		32'h00007B1A: begin
				q			<=			16'h0101;
		end
		32'h00007B1C: begin
				q			<=			16'h8067;
		end
		32'h00007B1E: begin
				q			<=			16'h0000;
		end
		32'h00007B20: begin
				q			<=			16'h2703;
		end
		32'h00007B22: begin
				q			<=			16'h0005;
		end
		32'h00007B24: begin
				q			<=			16'hA023;
		end
		32'h00007B26: begin
				q			<=			16'h00E7;
		end
		32'h00007B28: begin
				q			<=			16'h2823;
		end
		32'h00007B2A: begin
				q			<=			16'h0005;
		end
		32'h00007B2C: begin
				q			<=			16'h2623;
		end
		32'h00007B2E: begin
				q			<=			16'h0005;
		end
		32'h00007B30: begin
				q			<=			16'hF06F;
		end
		32'h00007B32: begin
				q			<=			16'hFD9F;
		end
		32'h00007B34: begin
				q			<=			16'h8063;
		end
		32'h00007B36: begin
				q			<=			16'h0205;
		end
		32'h00007B38: begin
				q			<=			16'hA783;
		end
		32'h00007B3A: begin
				q			<=			16'h0045;
		end
		32'h00007B3C: begin
				q			<=			16'h9713;
		end
		32'h00007B3E: begin
				q			<=			16'h0027;
		end
		32'h00007B40: begin
				q			<=			16'h2783;
		end
		32'h00007B42: begin
				q			<=			16'h04C5;
		end
		32'h00007B44: begin
				q			<=			16'h87B3;
		end
		32'h00007B46: begin
				q			<=			16'h00E7;
		end
		32'h00007B48: begin
				q			<=			16'hA703;
		end
		32'h00007B4A: begin
				q			<=			16'h0007;
		end
		32'h00007B4C: begin
				q			<=			16'hA023;
		end
		32'h00007B4E: begin
				q			<=			16'h00E5;
		end
		32'h00007B50: begin
				q			<=			16'hA023;
		end
		32'h00007B52: begin
				q			<=			16'h00B7;
		end
		32'h00007B54: begin
				q			<=			16'h8067;
		end
		32'h00007B56: begin
				q			<=			16'h0000;
		end
		32'h00007B58: begin
				q			<=			16'h0113;
		end
		32'h00007B5A: begin
				q			<=			16'hFD01;
		end
		32'h00007B5C: begin
				q			<=			16'h2E23;
		end
		32'h00007B5E: begin
				q			<=			16'h0131;
		end
		32'h00007B60: begin
				q			<=			16'h0993;
		end
		32'h00007B62: begin
				q			<=			16'h0005;
		end
		32'h00007B64: begin
				q			<=			16'h0537;
		end
		32'h00007B66: begin
				q			<=			16'h0001;
		end
		32'h00007B68: begin
				q			<=			16'h2423;
		end
		32'h00007B6A: begin
				q			<=			16'h0281;
		end
		32'h00007B6C: begin
				q			<=			16'h2223;
		end
		32'h00007B6E: begin
				q			<=			16'h0291;
		end
		32'h00007B70: begin
				q			<=			16'h8413;
		end
		32'h00007B72: begin
				q			<=			16'h0005;
		end
		32'h00007B74: begin
				q			<=			16'hA483;
		end
		32'h00007B76: begin
				q			<=			16'h0105;
		end
		32'h00007B78: begin
				q			<=			16'h2623;
		end
		32'h00007B7A: begin
				q			<=			16'h0211;
		end
		32'h00007B7C: begin
				q			<=			16'h2023;
		end
		32'h00007B7E: begin
				q			<=			16'h0321;
		end
		32'h00007B80: begin
				q			<=			16'h8593;
		end
		32'h00007B82: begin
				q			<=			16'h0145;
		end
		32'h00007B84: begin
				q			<=			16'h0813;
		end
		32'h00007B86: begin
				q			<=			16'h0000;
		end
		32'h00007B88: begin
				q			<=			16'h0513;
		end
		32'h00007B8A: begin
				q			<=			16'hFFF5;
		end
		32'h00007B8C: begin
				q			<=			16'hA783;
		end
		32'h00007B8E: begin
				q			<=			16'h0005;
		end
		32'h00007B90: begin
				q			<=			16'h8593;
		end
		32'h00007B92: begin
				q			<=			16'h0045;
		end
		32'h00007B94: begin
				q			<=			16'h0813;
		end
		32'h00007B96: begin
				q			<=			16'h0018;
		end
		32'h00007B98: begin
				q			<=			16'hF733;
		end
		32'h00007B9A: begin
				q			<=			16'h00A7;
		end
		32'h00007B9C: begin
				q			<=			16'h0733;
		end
		32'h00007B9E: begin
				q			<=			16'h02C7;
		end
		32'h00007BA0: begin
				q			<=			16'hD793;
		end
		32'h00007BA2: begin
				q			<=			16'h0107;
		end
		32'h00007BA4: begin
				q			<=			16'h87B3;
		end
		32'h00007BA6: begin
				q			<=			16'h02C7;
		end
		32'h00007BA8: begin
				q			<=			16'h0733;
		end
		32'h00007BAA: begin
				q			<=			16'h00D7;
		end
		32'h00007BAC: begin
				q			<=			16'h5693;
		end
		32'h00007BAE: begin
				q			<=			16'h0107;
		end
		32'h00007BB0: begin
				q			<=			16'h7733;
		end
		32'h00007BB2: begin
				q			<=			16'h00A7;
		end
		32'h00007BB4: begin
				q			<=			16'h87B3;
		end
		32'h00007BB6: begin
				q			<=			16'h00D7;
		end
		32'h00007BB8: begin
				q			<=			16'hD693;
		end
		32'h00007BBA: begin
				q			<=			16'h0107;
		end
		32'h00007BBC: begin
				q			<=			16'h9793;
		end
		32'h00007BBE: begin
				q			<=			16'h0107;
		end
		32'h00007BC0: begin
				q			<=			16'h87B3;
		end
		32'h00007BC2: begin
				q			<=			16'h00E7;
		end
		32'h00007BC4: begin
				q			<=			16'hAE23;
		end
		32'h00007BC6: begin
				q			<=			16'hFEF5;
		end
		32'h00007BC8: begin
				q			<=			16'h42E3;
		end
		32'h00007BCA: begin
				q			<=			16'hFC98;
		end
		32'h00007BCC: begin
				q			<=			16'h8663;
		end
		32'h00007BCE: begin
				q			<=			16'h0606;
		end
		32'h00007BD0: begin
				q			<=			16'h2783;
		end
		32'h00007BD2: begin
				q			<=			16'h0084;
		end
		32'h00007BD4: begin
				q			<=			16'hC663;
		end
		32'h00007BD6: begin
				q			<=			16'h04F4;
		end
		32'h00007BD8: begin
				q			<=			16'h2583;
		end
		32'h00007BDA: begin
				q			<=			16'h0044;
		end
		32'h00007BDC: begin
				q			<=			16'h8513;
		end
		32'h00007BDE: begin
				q			<=			16'h0009;
		end
		32'h00007BE0: begin
				q			<=			16'h2623;
		end
		32'h00007BE2: begin
				q			<=			16'h00D1;
		end
		32'h00007BE4: begin
				q			<=			16'h8593;
		end
		32'h00007BE6: begin
				q			<=			16'h0015;
		end
		32'h00007BE8: begin
				q			<=			16'hF0EF;
		end
		32'h00007BEA: begin
				q			<=			16'hEA5F;
		end
		32'h00007BEC: begin
				q			<=			16'h2603;
		end
		32'h00007BEE: begin
				q			<=			16'h0104;
		end
		32'h00007BF0: begin
				q			<=			16'h0593;
		end
		32'h00007BF2: begin
				q			<=			16'h00C4;
		end
		32'h00007BF4: begin
				q			<=			16'h0913;
		end
		32'h00007BF6: begin
				q			<=			16'h0005;
		end
		32'h00007BF8: begin
				q			<=			16'h0613;
		end
		32'h00007BFA: begin
				q			<=			16'h0026;
		end
		32'h00007BFC: begin
				q			<=			16'h1613;
		end
		32'h00007BFE: begin
				q			<=			16'h0026;
		end
		32'h00007C00: begin
				q			<=			16'h0513;
		end
		32'h00007C02: begin
				q			<=			16'h00C5;
		end
		32'h00007C04: begin
				q			<=			16'hA0EF;
		end
		32'h00007C06: begin
				q			<=			16'hEF5F;
		end
		32'h00007C08: begin
				q			<=			16'h0593;
		end
		32'h00007C0A: begin
				q			<=			16'h0004;
		end
		32'h00007C0C: begin
				q			<=			16'h8513;
		end
		32'h00007C0E: begin
				q			<=			16'h0009;
		end
		32'h00007C10: begin
				q			<=			16'h0097;
		end
		32'h00007C12: begin
				q			<=			16'h0000;
		end
		32'h00007C14: begin
				q			<=			16'h80E7;
		end
		32'h00007C16: begin
				q			<=			16'hF240;
		end
		32'h00007C18: begin
				q			<=			16'h2683;
		end
		32'h00007C1A: begin
				q			<=			16'h00C1;
		end
		32'h00007C1C: begin
				q			<=			16'h0413;
		end
		32'h00007C1E: begin
				q			<=			16'h0009;
		end
		32'h00007C20: begin
				q			<=			16'h8793;
		end
		32'h00007C22: begin
				q			<=			16'h0044;
		end
		32'h00007C24: begin
				q			<=			16'h9793;
		end
		32'h00007C26: begin
				q			<=			16'h0027;
		end
		32'h00007C28: begin
				q			<=			16'h07B3;
		end
		32'h00007C2A: begin
				q			<=			16'h00F4;
		end
		32'h00007C2C: begin
				q			<=			16'hA223;
		end
		32'h00007C2E: begin
				q			<=			16'h00D7;
		end
		32'h00007C30: begin
				q			<=			16'h8493;
		end
		32'h00007C32: begin
				q			<=			16'h0014;
		end
		32'h00007C34: begin
				q			<=			16'h2823;
		end
		32'h00007C36: begin
				q			<=			16'h0094;
		end
		32'h00007C38: begin
				q			<=			16'h0513;
		end
		32'h00007C3A: begin
				q			<=			16'h0004;
		end
		32'h00007C3C: begin
				q			<=			16'h2083;
		end
		32'h00007C3E: begin
				q			<=			16'h02C1;
		end
		32'h00007C40: begin
				q			<=			16'h2403;
		end
		32'h00007C42: begin
				q			<=			16'h0281;
		end
		32'h00007C44: begin
				q			<=			16'h2483;
		end
		32'h00007C46: begin
				q			<=			16'h0241;
		end
		32'h00007C48: begin
				q			<=			16'h2903;
		end
		32'h00007C4A: begin
				q			<=			16'h0201;
		end
		32'h00007C4C: begin
				q			<=			16'h2983;
		end
		32'h00007C4E: begin
				q			<=			16'h01C1;
		end
		32'h00007C50: begin
				q			<=			16'h0113;
		end
		32'h00007C52: begin
				q			<=			16'h0301;
		end
		32'h00007C54: begin
				q			<=			16'h8067;
		end
		32'h00007C56: begin
				q			<=			16'h0000;
		end
		32'h00007C58: begin
				q			<=			16'h0113;
		end
		32'h00007C5A: begin
				q			<=			16'hFD01;
		end
		32'h00007C5C: begin
				q			<=			16'h8793;
		end
		32'h00007C5E: begin
				q			<=			16'h0086;
		end
		32'h00007C60: begin
				q			<=			16'h2C23;
		end
		32'h00007C62: begin
				q			<=			16'h0141;
		end
		32'h00007C64: begin
				q			<=			16'h8A13;
		end
		32'h00007C66: begin
				q			<=			16'h0006;
		end
		32'h00007C68: begin
				q			<=			16'h0693;
		end
		32'h00007C6A: begin
				q			<=			16'h0090;
		end
		32'h00007C6C: begin
				q			<=			16'h2423;
		end
		32'h00007C6E: begin
				q			<=			16'h0281;
		end
		32'h00007C70: begin
				q			<=			16'h2223;
		end
		32'h00007C72: begin
				q			<=			16'h0291;
		end
		32'h00007C74: begin
				q			<=			16'h2E23;
		end
		32'h00007C76: begin
				q			<=			16'h0131;
		end
		32'h00007C78: begin
				q			<=			16'h8413;
		end
		32'h00007C7A: begin
				q			<=			16'h0005;
		end
		32'h00007C7C: begin
				q			<=			16'hC7B3;
		end
		32'h00007C7E: begin
				q			<=			16'h02D7;
		end
		32'h00007C80: begin
				q			<=			16'h2623;
		end
		32'h00007C82: begin
				q			<=			16'h0211;
		end
		32'h00007C84: begin
				q			<=			16'h2023;
		end
		32'h00007C86: begin
				q			<=			16'h0321;
		end
		32'h00007C88: begin
				q			<=			16'h2A23;
		end
		32'h00007C8A: begin
				q			<=			16'h0151;
		end
		32'h00007C8C: begin
				q			<=			16'h0993;
		end
		32'h00007C8E: begin
				q			<=			16'h0005;
		end
		32'h00007C90: begin
				q			<=			16'h0493;
		end
		32'h00007C92: begin
				q			<=			16'h0006;
		end
		32'h00007C94: begin
				q			<=			16'h0693;
		end
		32'h00007C96: begin
				q			<=			16'h0010;
		end
		32'h00007C98: begin
				q			<=			16'h0593;
		end
		32'h00007C9A: begin
				q			<=			16'h0000;
		end
		32'h00007C9C: begin
				q			<=			16'hCA63;
		end
		32'h00007C9E: begin
				q			<=			16'h08F6;
		end
		32'h00007CA0: begin
				q			<=			16'h8513;
		end
		32'h00007CA2: begin
				q			<=			16'h0009;
		end
		32'h00007CA4: begin
				q			<=			16'h2623;
		end
		32'h00007CA6: begin
				q			<=			16'h00E1;
		end
		32'h00007CA8: begin
				q			<=			16'h0097;
		end
		32'h00007CAA: begin
				q			<=			16'h0000;
		end
		32'h00007CAC: begin
				q			<=			16'h80E7;
		end
		32'h00007CAE: begin
				q			<=			16'hDE40;
		end
		32'h00007CB0: begin
				q			<=			16'h2703;
		end
		32'h00007CB2: begin
				q			<=			16'h00C1;
		end
		32'h00007CB4: begin
				q			<=			16'h0793;
		end
		32'h00007CB6: begin
				q			<=			16'h0010;
		end
		32'h00007CB8: begin
				q			<=			16'h2823;
		end
		32'h00007CBA: begin
				q			<=			16'h00F5;
		end
		32'h00007CBC: begin
				q			<=			16'h2A23;
		end
		32'h00007CBE: begin
				q			<=			16'h00E5;
		end
		32'h00007CC0: begin
				q			<=			16'h0793;
		end
		32'h00007CC2: begin
				q			<=			16'h0090;
		end
		32'h00007CC4: begin
				q			<=			16'hDC63;
		end
		32'h00007CC6: begin
				q			<=			16'h0697;
		end
		32'h00007CC8: begin
				q			<=			16'h0A93;
		end
		32'h00007CCA: begin
				q			<=			16'h0094;
		end
		32'h00007CCC: begin
				q			<=			16'h8913;
		end
		32'h00007CCE: begin
				q			<=			16'h000A;
		end
		32'h00007CD0: begin
				q			<=			16'h0433;
		end
		32'h00007CD2: begin
				q			<=			16'h0094;
		end
		32'h00007CD4: begin
				q			<=			16'h0913;
		end
		32'h00007CD6: begin
				q			<=			16'h0019;
		end
		32'h00007CD8: begin
				q			<=			16'h4683;
		end
		32'h00007CDA: begin
				q			<=			16'hFFF9;
		end
		32'h00007CDC: begin
				q			<=			16'h0593;
		end
		32'h00007CDE: begin
				q			<=			16'h0005;
		end
		32'h00007CE0: begin
				q			<=			16'h0613;
		end
		32'h00007CE2: begin
				q			<=			16'h00A0;
		end
		32'h00007CE4: begin
				q			<=			16'h8693;
		end
		32'h00007CE6: begin
				q			<=			16'hFD06;
		end
		32'h00007CE8: begin
				q			<=			16'h8513;
		end
		32'h00007CEA: begin
				q			<=			16'h0009;
		end
		32'h00007CEC: begin
				q			<=			16'h0097;
		end
		32'h00007CEE: begin
				q			<=			16'h0000;
		end
		32'h00007CF0: begin
				q			<=			16'h80E7;
		end
		32'h00007CF2: begin
				q			<=			16'hE6C0;
		end
		32'h00007CF4: begin
				q			<=			16'h10E3;
		end
		32'h00007CF6: begin
				q			<=			16'hFE89;
		end
		32'h00007CF8: begin
				q			<=			16'h8413;
		end
		32'h00007CFA: begin
				q			<=			16'hFF84;
		end
		32'h00007CFC: begin
				q			<=			16'h8433;
		end
		32'h00007CFE: begin
				q			<=			16'h008A;
		end
		32'h00007D00: begin
				q			<=			16'h84B3;
		end
		32'h00007D02: begin
				q			<=			16'h4084;
		end
		32'h00007D04: begin
				q			<=			16'h07B3;
		end
		32'h00007D06: begin
				q			<=			16'h0094;
		end
		32'h00007D08: begin
				q			<=			16'hC063;
		end
		32'h00007D0A: begin
				q			<=			16'h0547;
		end
		32'h00007D0C: begin
				q			<=			16'h2083;
		end
		32'h00007D0E: begin
				q			<=			16'h02C1;
		end
		32'h00007D10: begin
				q			<=			16'h2403;
		end
		32'h00007D12: begin
				q			<=			16'h0281;
		end
		32'h00007D14: begin
				q			<=			16'h2483;
		end
		32'h00007D16: begin
				q			<=			16'h0241;
		end
		32'h00007D18: begin
				q			<=			16'h2903;
		end
		32'h00007D1A: begin
				q			<=			16'h0201;
		end
		32'h00007D1C: begin
				q			<=			16'h2983;
		end
		32'h00007D1E: begin
				q			<=			16'h01C1;
		end
		32'h00007D20: begin
				q			<=			16'h2A03;
		end
		32'h00007D22: begin
				q			<=			16'h0181;
		end
		32'h00007D24: begin
				q			<=			16'h2A83;
		end
		32'h00007D26: begin
				q			<=			16'h0141;
		end
		32'h00007D28: begin
				q			<=			16'h0113;
		end
		32'h00007D2A: begin
				q			<=			16'h0301;
		end
		32'h00007D2C: begin
				q			<=			16'h8067;
		end
		32'h00007D2E: begin
				q			<=			16'h0000;
		end
		32'h00007D30: begin
				q			<=			16'h9693;
		end
		32'h00007D32: begin
				q			<=			16'h0016;
		end
		32'h00007D34: begin
				q			<=			16'h8593;
		end
		32'h00007D36: begin
				q			<=			16'h0015;
		end
		32'h00007D38: begin
				q			<=			16'hF06F;
		end
		32'h00007D3A: begin
				q			<=			16'hF65F;
		end
		32'h00007D3C: begin
				q			<=			16'h0413;
		end
		32'h00007D3E: begin
				q			<=			16'h00A4;
		end
		32'h00007D40: begin
				q			<=			16'h0493;
		end
		32'h00007D42: begin
				q			<=			16'h0090;
		end
		32'h00007D44: begin
				q			<=			16'hF06F;
		end
		32'h00007D46: begin
				q			<=			16'hFBDF;
		end
		32'h00007D48: begin
				q			<=			16'h0413;
		end
		32'h00007D4A: begin
				q			<=			16'h0014;
		end
		32'h00007D4C: begin
				q			<=			16'h4683;
		end
		32'h00007D4E: begin
				q			<=			16'hFFF4;
		end
		32'h00007D50: begin
				q			<=			16'h0593;
		end
		32'h00007D52: begin
				q			<=			16'h0005;
		end
		32'h00007D54: begin
				q			<=			16'h0613;
		end
		32'h00007D56: begin
				q			<=			16'h00A0;
		end
		32'h00007D58: begin
				q			<=			16'h8693;
		end
		32'h00007D5A: begin
				q			<=			16'hFD06;
		end
		32'h00007D5C: begin
				q			<=			16'h8513;
		end
		32'h00007D5E: begin
				q			<=			16'h0009;
		end
		32'h00007D60: begin
				q			<=			16'h0097;
		end
		32'h00007D62: begin
				q			<=			16'h0000;
		end
		32'h00007D64: begin
				q			<=			16'h80E7;
		end
		32'h00007D66: begin
				q			<=			16'hDF80;
		end
		32'h00007D68: begin
				q			<=			16'hF06F;
		end
		32'h00007D6A: begin
				q			<=			16'hF9DF;
		end
		32'h00007D6C: begin
				q			<=			16'h0737;
		end
		32'h00007D6E: begin
				q			<=			16'hFFFF;
		end
		32'h00007D70: begin
				q			<=			16'h7733;
		end
		32'h00007D72: begin
				q			<=			16'h00E5;
		end
		32'h00007D74: begin
				q			<=			16'h0793;
		end
		32'h00007D76: begin
				q			<=			16'h0005;
		end
		32'h00007D78: begin
				q			<=			16'h0513;
		end
		32'h00007D7A: begin
				q			<=			16'h0000;
		end
		32'h00007D7C: begin
				q			<=			16'h1663;
		end
		32'h00007D7E: begin
				q			<=			16'h0007;
		end
		32'h00007D80: begin
				q			<=			16'h9793;
		end
		32'h00007D82: begin
				q			<=			16'h0107;
		end
		32'h00007D84: begin
				q			<=			16'h0513;
		end
		32'h00007D86: begin
				q			<=			16'h0100;
		end
		32'h00007D88: begin
				q			<=			16'h0737;
		end
		32'h00007D8A: begin
				q			<=			16'hFF00;
		end
		32'h00007D8C: begin
				q			<=			16'hF733;
		end
		32'h00007D8E: begin
				q			<=			16'h00E7;
		end
		32'h00007D90: begin
				q			<=			16'h1663;
		end
		32'h00007D92: begin
				q			<=			16'h0007;
		end
		32'h00007D94: begin
				q			<=			16'h0513;
		end
		32'h00007D96: begin
				q			<=			16'h0085;
		end
		32'h00007D98: begin
				q			<=			16'h9793;
		end
		32'h00007D9A: begin
				q			<=			16'h0087;
		end
		32'h00007D9C: begin
				q			<=			16'h0737;
		end
		32'h00007D9E: begin
				q			<=			16'hF000;
		end
		32'h00007DA0: begin
				q			<=			16'hF733;
		end
		32'h00007DA2: begin
				q			<=			16'h00E7;
		end
		32'h00007DA4: begin
				q			<=			16'h1663;
		end
		32'h00007DA6: begin
				q			<=			16'h0007;
		end
		32'h00007DA8: begin
				q			<=			16'h0513;
		end
		32'h00007DAA: begin
				q			<=			16'h0045;
		end
		32'h00007DAC: begin
				q			<=			16'h9793;
		end
		32'h00007DAE: begin
				q			<=			16'h0047;
		end
		32'h00007DB0: begin
				q			<=			16'h0737;
		end
		32'h00007DB2: begin
				q			<=			16'hC000;
		end
		32'h00007DB4: begin
				q			<=			16'hF733;
		end
		32'h00007DB6: begin
				q			<=			16'h00E7;
		end
		32'h00007DB8: begin
				q			<=			16'h1663;
		end
		32'h00007DBA: begin
				q			<=			16'h0007;
		end
		32'h00007DBC: begin
				q			<=			16'h0513;
		end
		32'h00007DBE: begin
				q			<=			16'h0025;
		end
		32'h00007DC0: begin
				q			<=			16'h9793;
		end
		32'h00007DC2: begin
				q			<=			16'h0027;
		end
		32'h00007DC4: begin
				q			<=			16'hCC63;
		end
		32'h00007DC6: begin
				q			<=			16'h0007;
		end
		32'h00007DC8: begin
				q			<=			16'h9713;
		end
		32'h00007DCA: begin
				q			<=			16'h0017;
		end
		32'h00007DCC: begin
				q			<=			16'h5663;
		end
		32'h00007DCE: begin
				q			<=			16'h0007;
		end
		32'h00007DD0: begin
				q			<=			16'h0513;
		end
		32'h00007DD2: begin
				q			<=			16'h0015;
		end
		32'h00007DD4: begin
				q			<=			16'h8067;
		end
		32'h00007DD6: begin
				q			<=			16'h0000;
		end
		32'h00007DD8: begin
				q			<=			16'h0513;
		end
		32'h00007DDA: begin
				q			<=			16'h0200;
		end
		32'h00007DDC: begin
				q			<=			16'h8067;
		end
		32'h00007DDE: begin
				q			<=			16'h0000;
		end
		32'h00007DE0: begin
				q			<=			16'h2783;
		end
		32'h00007DE2: begin
				q			<=			16'h0005;
		end
		32'h00007DE4: begin
				q			<=			16'hF713;
		end
		32'h00007DE6: begin
				q			<=			16'h0077;
		end
		32'h00007DE8: begin
				q			<=			16'h0E63;
		end
		32'h00007DEA: begin
				q			<=			16'h0207;
		end
		32'h00007DEC: begin
				q			<=			16'hF693;
		end
		32'h00007DEE: begin
				q			<=			16'h0017;
		end
		32'h00007DF0: begin
				q			<=			16'h0713;
		end
		32'h00007DF2: begin
				q			<=			16'h0000;
		end
		32'h00007DF4: begin
				q			<=			16'h9C63;
		end
		32'h00007DF6: begin
				q			<=			16'h0006;
		end
		32'h00007DF8: begin
				q			<=			16'hF713;
		end
		32'h00007DFA: begin
				q			<=			16'h0027;
		end
		32'h00007DFC: begin
				q			<=			16'h0C63;
		end
		32'h00007DFE: begin
				q			<=			16'h0007;
		end
		32'h00007E00: begin
				q			<=			16'hD793;
		end
		32'h00007E02: begin
				q			<=			16'h0017;
		end
		32'h00007E04: begin
				q			<=			16'h2023;
		end
		32'h00007E06: begin
				q			<=			16'h00F5;
		end
		32'h00007E08: begin
				q			<=			16'h0713;
		end
		32'h00007E0A: begin
				q			<=			16'h0010;
		end
		32'h00007E0C: begin
				q			<=			16'h0513;
		end
		32'h00007E0E: begin
				q			<=			16'h0007;
		end
		32'h00007E10: begin
				q			<=			16'h8067;
		end
		32'h00007E12: begin
				q			<=			16'h0000;
		end
		32'h00007E14: begin
				q			<=			16'hD793;
		end
		32'h00007E16: begin
				q			<=			16'h0027;
		end
		32'h00007E18: begin
				q			<=			16'h2023;
		end
		32'h00007E1A: begin
				q			<=			16'h00F5;
		end
		32'h00007E1C: begin
				q			<=			16'h0713;
		end
		32'h00007E1E: begin
				q			<=			16'h0020;
		end
		32'h00007E20: begin
				q			<=			16'hF06F;
		end
		32'h00007E22: begin
				q			<=			16'hFEDF;
		end
		32'h00007E24: begin
				q			<=			16'h9693;
		end
		32'h00007E26: begin
				q			<=			16'h0107;
		end
		32'h00007E28: begin
				q			<=			16'hD693;
		end
		32'h00007E2A: begin
				q			<=			16'h0106;
		end
		32'h00007E2C: begin
				q			<=			16'h0713;
		end
		32'h00007E2E: begin
				q			<=			16'h0000;
		end
		32'h00007E30: begin
				q			<=			16'h9663;
		end
		32'h00007E32: begin
				q			<=			16'h0006;
		end
		32'h00007E34: begin
				q			<=			16'hD793;
		end
		32'h00007E36: begin
				q			<=			16'h0107;
		end
		32'h00007E38: begin
				q			<=			16'h0713;
		end
		32'h00007E3A: begin
				q			<=			16'h0100;
		end
		32'h00007E3C: begin
				q			<=			16'hF693;
		end
		32'h00007E3E: begin
				q			<=			16'h0FF7;
		end
		32'h00007E40: begin
				q			<=			16'h9663;
		end
		32'h00007E42: begin
				q			<=			16'h0006;
		end
		32'h00007E44: begin
				q			<=			16'h0713;
		end
		32'h00007E46: begin
				q			<=			16'h0087;
		end
		32'h00007E48: begin
				q			<=			16'hD793;
		end
		32'h00007E4A: begin
				q			<=			16'h0087;
		end
		32'h00007E4C: begin
				q			<=			16'hF693;
		end
		32'h00007E4E: begin
				q			<=			16'h00F7;
		end
		32'h00007E50: begin
				q			<=			16'h9663;
		end
		32'h00007E52: begin
				q			<=			16'h0006;
		end
		32'h00007E54: begin
				q			<=			16'h0713;
		end
		32'h00007E56: begin
				q			<=			16'h0047;
		end
		32'h00007E58: begin
				q			<=			16'hD793;
		end
		32'h00007E5A: begin
				q			<=			16'h0047;
		end
		32'h00007E5C: begin
				q			<=			16'hF693;
		end
		32'h00007E5E: begin
				q			<=			16'h0037;
		end
		32'h00007E60: begin
				q			<=			16'h9663;
		end
		32'h00007E62: begin
				q			<=			16'h0006;
		end
		32'h00007E64: begin
				q			<=			16'h0713;
		end
		32'h00007E66: begin
				q			<=			16'h0027;
		end
		32'h00007E68: begin
				q			<=			16'hD793;
		end
		32'h00007E6A: begin
				q			<=			16'h0027;
		end
		32'h00007E6C: begin
				q			<=			16'hF693;
		end
		32'h00007E6E: begin
				q			<=			16'h0017;
		end
		32'h00007E70: begin
				q			<=			16'h9863;
		end
		32'h00007E72: begin
				q			<=			16'h0006;
		end
		32'h00007E74: begin
				q			<=			16'hD793;
		end
		32'h00007E76: begin
				q			<=			16'h0017;
		end
		32'h00007E78: begin
				q			<=			16'h8863;
		end
		32'h00007E7A: begin
				q			<=			16'h0007;
		end
		32'h00007E7C: begin
				q			<=			16'h0713;
		end
		32'h00007E7E: begin
				q			<=			16'h0017;
		end
		32'h00007E80: begin
				q			<=			16'h2023;
		end
		32'h00007E82: begin
				q			<=			16'h00F5;
		end
		32'h00007E84: begin
				q			<=			16'hF06F;
		end
		32'h00007E86: begin
				q			<=			16'hF89F;
		end
		32'h00007E88: begin
				q			<=			16'h0713;
		end
		32'h00007E8A: begin
				q			<=			16'h0200;
		end
		32'h00007E8C: begin
				q			<=			16'hF06F;
		end
		32'h00007E8E: begin
				q			<=			16'hF81F;
		end
		32'h00007E90: begin
				q			<=			16'h0113;
		end
		32'h00007E92: begin
				q			<=			16'hFF01;
		end
		32'h00007E94: begin
				q			<=			16'h2423;
		end
		32'h00007E96: begin
				q			<=			16'h0081;
		end
		32'h00007E98: begin
				q			<=			16'h8413;
		end
		32'h00007E9A: begin
				q			<=			16'h0005;
		end
		32'h00007E9C: begin
				q			<=			16'h0593;
		end
		32'h00007E9E: begin
				q			<=			16'h0010;
		end
		32'h00007EA0: begin
				q			<=			16'h2623;
		end
		32'h00007EA2: begin
				q			<=			16'h0011;
		end
		32'h00007EA4: begin
				q			<=			16'hF0EF;
		end
		32'h00007EA6: begin
				q			<=			16'hBE9F;
		end
		32'h00007EA8: begin
				q			<=			16'h2A23;
		end
		32'h00007EAA: begin
				q			<=			16'h0085;
		end
		32'h00007EAC: begin
				q			<=			16'h2083;
		end
		32'h00007EAE: begin
				q			<=			16'h00C1;
		end
		32'h00007EB0: begin
				q			<=			16'h2403;
		end
		32'h00007EB2: begin
				q			<=			16'h0081;
		end
		32'h00007EB4: begin
				q			<=			16'h0713;
		end
		32'h00007EB6: begin
				q			<=			16'h0010;
		end
		32'h00007EB8: begin
				q			<=			16'h2823;
		end
		32'h00007EBA: begin
				q			<=			16'h00E5;
		end
		32'h00007EBC: begin
				q			<=			16'h0113;
		end
		32'h00007EBE: begin
				q			<=			16'h0101;
		end
		32'h00007EC0: begin
				q			<=			16'h8067;
		end
		32'h00007EC2: begin
				q			<=			16'h0000;
		end
		32'h00007EC4: begin
				q			<=			16'hA703;
		end
		32'h00007EC6: begin
				q			<=			16'h0105;
		end
		32'h00007EC8: begin
				q			<=			16'h2783;
		end
		32'h00007ECA: begin
				q			<=			16'h0106;
		end
		32'h00007ECC: begin
				q			<=			16'h0113;
		end
		32'h00007ECE: begin
				q			<=			16'hFD01;
		end
		32'h00007ED0: begin
				q			<=			16'h2223;
		end
		32'h00007ED2: begin
				q			<=			16'h0291;
		end
		32'h00007ED4: begin
				q			<=			16'h2623;
		end
		32'h00007ED6: begin
				q			<=			16'h0211;
		end
		32'h00007ED8: begin
				q			<=			16'h2423;
		end
		32'h00007EDA: begin
				q			<=			16'h0281;
		end
		32'h00007EDC: begin
				q			<=			16'h2023;
		end
		32'h00007EDE: begin
				q			<=			16'h0321;
		end
		32'h00007EE0: begin
				q			<=			16'h2E23;
		end
		32'h00007EE2: begin
				q			<=			16'h0131;
		end
		32'h00007EE4: begin
				q			<=			16'h8493;
		end
		32'h00007EE6: begin
				q			<=			16'h0005;
		end
		32'h00007EE8: begin
				q			<=			16'h5663;
		end
		32'h00007EEA: begin
				q			<=			16'h00F7;
		end
		32'h00007EEC: begin
				q			<=			16'h0493;
		end
		32'h00007EEE: begin
				q			<=			16'h0006;
		end
		32'h00007EF0: begin
				q			<=			16'h8613;
		end
		32'h00007EF2: begin
				q			<=			16'h0005;
		end
		32'h00007EF4: begin
				q			<=			16'hA983;
		end
		32'h00007EF6: begin
				q			<=			16'h0104;
		end
		32'h00007EF8: begin
				q			<=			16'h2903;
		end
		32'h00007EFA: begin
				q			<=			16'h0106;
		end
		32'h00007EFC: begin
				q			<=			16'hA783;
		end
		32'h00007EFE: begin
				q			<=			16'h0084;
		end
		32'h00007F00: begin
				q			<=			16'hA583;
		end
		32'h00007F02: begin
				q			<=			16'h0044;
		end
		32'h00007F04: begin
				q			<=			16'h8433;
		end
		32'h00007F06: begin
				q			<=			16'h0129;
		end
		32'h00007F08: begin
				q			<=			16'hD463;
		end
		32'h00007F0A: begin
				q			<=			16'h0087;
		end
		32'h00007F0C: begin
				q			<=			16'h8593;
		end
		32'h00007F0E: begin
				q			<=			16'h0015;
		end
		32'h00007F10: begin
				q			<=			16'h2623;
		end
		32'h00007F12: begin
				q			<=			16'h00C1;
		end
		32'h00007F14: begin
				q			<=			16'h0097;
		end
		32'h00007F16: begin
				q			<=			16'h0000;
		end
		32'h00007F18: begin
				q			<=			16'h80E7;
		end
		32'h00007F1A: begin
				q			<=			16'hB780;
		end
		32'h00007F1C: begin
				q			<=			16'h2603;
		end
		32'h00007F1E: begin
				q			<=			16'h00C1;
		end
		32'h00007F20: begin
				q			<=			16'h0813;
		end
		32'h00007F22: begin
				q			<=			16'h0145;
		end
		32'h00007F24: begin
				q			<=			16'h1313;
		end
		32'h00007F26: begin
				q			<=			16'h0024;
		end
		32'h00007F28: begin
				q			<=			16'h0333;
		end
		32'h00007F2A: begin
				q			<=			16'h0068;
		end
		32'h00007F2C: begin
				q			<=			16'h0793;
		end
		32'h00007F2E: begin
				q			<=			16'h0008;
		end
		32'h00007F30: begin
				q			<=			16'hEC63;
		end
		32'h00007F32: begin
				q			<=			16'h0467;
		end
		32'h00007F34: begin
				q			<=			16'h8593;
		end
		32'h00007F36: begin
				q			<=			16'h0144;
		end
		32'h00007F38: begin
				q			<=			16'h9893;
		end
		32'h00007F3A: begin
				q			<=			16'h0029;
		end
		32'h00007F3C: begin
				q			<=			16'h0613;
		end
		32'h00007F3E: begin
				q			<=			16'h0146;
		end
		32'h00007F40: begin
				q			<=			16'h1E13;
		end
		32'h00007F42: begin
				q			<=			16'h0029;
		end
		32'h00007F44: begin
				q			<=			16'h06B7;
		end
		32'h00007F46: begin
				q			<=			16'h0001;
		end
		32'h00007F48: begin
				q			<=			16'h88B3;
		end
		32'h00007F4A: begin
				q			<=			16'h0115;
		end
		32'h00007F4C: begin
				q			<=			16'h0E33;
		end
		32'h00007F4E: begin
				q			<=			16'h01C6;
		end
		32'h00007F50: begin
				q			<=			16'h8693;
		end
		32'h00007F52: begin
				q			<=			16'hFFF6;
		end
		32'h00007F54: begin
				q			<=			16'h6063;
		end
		32'h00007F56: begin
				q			<=			16'h05C6;
		end
		32'h00007F58: begin
				q			<=			16'h5863;
		end
		32'h00007F5A: begin
				q			<=			16'h0080;
		end
		32'h00007F5C: begin
				q			<=			16'h0313;
		end
		32'h00007F5E: begin
				q			<=			16'hFFC3;
		end
		32'h00007F60: begin
				q			<=			16'h2783;
		end
		32'h00007F62: begin
				q			<=			16'h0003;
		end
		32'h00007F64: begin
				q			<=			16'h8E63;
		end
		32'h00007F66: begin
				q			<=			16'h1007;
		end
		32'h00007F68: begin
				q			<=			16'h2823;
		end
		32'h00007F6A: begin
				q			<=			16'h0085;
		end
		32'h00007F6C: begin
				q			<=			16'h2083;
		end
		32'h00007F6E: begin
				q			<=			16'h02C1;
		end
		32'h00007F70: begin
				q			<=			16'h2403;
		end
		32'h00007F72: begin
				q			<=			16'h0281;
		end
		32'h00007F74: begin
				q			<=			16'h2483;
		end
		32'h00007F76: begin
				q			<=			16'h0241;
		end
		32'h00007F78: begin
				q			<=			16'h2903;
		end
		32'h00007F7A: begin
				q			<=			16'h0201;
		end
		32'h00007F7C: begin
				q			<=			16'h2983;
		end
		32'h00007F7E: begin
				q			<=			16'h01C1;
		end
		32'h00007F80: begin
				q			<=			16'h0113;
		end
		32'h00007F82: begin
				q			<=			16'h0301;
		end
		32'h00007F84: begin
				q			<=			16'h8067;
		end
		32'h00007F86: begin
				q			<=			16'h0000;
		end
		32'h00007F88: begin
				q			<=			16'hA023;
		end
		32'h00007F8A: begin
				q			<=			16'h0007;
		end
		32'h00007F8C: begin
				q			<=			16'h8793;
		end
		32'h00007F8E: begin
				q			<=			16'h0047;
		end
		32'h00007F90: begin
				q			<=			16'hF06F;
		end
		32'h00007F92: begin
				q			<=			16'hFA1F;
		end
		32'h00007F94: begin
				q			<=			16'h2F83;
		end
		32'h00007F96: begin
				q			<=			16'h0006;
		end
		32'h00007F98: begin
				q			<=			16'hFFB3;
		end
		32'h00007F9A: begin
				q			<=			16'h00DF;
		end
		32'h00007F9C: begin
				q			<=			16'h8463;
		end
		32'h00007F9E: begin
				q			<=			16'h060F;
		end
		32'h00007FA0: begin
				q			<=			16'h0F13;
		end
		32'h00007FA2: begin
				q			<=			16'h0008;
		end
		32'h00007FA4: begin
				q			<=			16'h8293;
		end
		32'h00007FA6: begin
				q			<=			16'h0005;
		end
		32'h00007FA8: begin
				q			<=			16'h0493;
		end
		32'h00007FAA: begin
				q			<=			16'h0000;
		end
		32'h00007FAC: begin
				q			<=			16'hA703;
		end
		32'h00007FAE: begin
				q			<=			16'h0002;
		end
		32'h00007FB0: begin
				q			<=			16'h2383;
		end
		32'h00007FB2: begin
				q			<=			16'h000F;
		end
		32'h00007FB4: begin
				q			<=			16'h0F13;
		end
		32'h00007FB6: begin
				q			<=			16'h004F;
		end
		32'h00007FB8: begin
				q			<=			16'h7EB3;
		end
		32'h00007FBA: begin
				q			<=			16'h00D7;
		end
		32'h00007FBC: begin
				q			<=			16'h8EB3;
		end
		32'h00007FBE: begin
				q			<=			16'h03FE;
		end
		32'h00007FC0: begin
				q			<=			16'hF7B3;
		end
		32'h00007FC2: begin
				q			<=			16'h00D3;
		end
		32'h00007FC4: begin
				q			<=			16'hD393;
		end
		32'h00007FC6: begin
				q			<=			16'h0103;
		end
		32'h00007FC8: begin
				q			<=			16'h8293;
		end
		32'h00007FCA: begin
				q			<=			16'h0042;
		end
		32'h00007FCC: begin
				q			<=			16'h8EB3;
		end
		32'h00007FCE: begin
				q			<=			16'h00FE;
		end
		32'h00007FD0: begin
				q			<=			16'h5793;
		end
		32'h00007FD2: begin
				q			<=			16'h0107;
		end
		32'h00007FD4: begin
				q			<=			16'h87B3;
		end
		32'h00007FD6: begin
				q			<=			16'h03F7;
		end
		32'h00007FD8: begin
				q			<=			16'h8EB3;
		end
		32'h00007FDA: begin
				q			<=			16'h009E;
		end
		32'h00007FDC: begin
				q			<=			16'hD713;
		end
		32'h00007FDE: begin
				q			<=			16'h010E;
		end
		32'h00007FE0: begin
				q			<=			16'hFEB3;
		end
		32'h00007FE2: begin
				q			<=			16'h00DE;
		end
		32'h00007FE4: begin
				q			<=			16'h87B3;
		end
		32'h00007FE6: begin
				q			<=			16'h0077;
		end
		32'h00007FE8: begin
				q			<=			16'h87B3;
		end
		32'h00007FEA: begin
				q			<=			16'h00E7;
		end
		32'h00007FEC: begin
				q			<=			16'hD493;
		end
		32'h00007FEE: begin
				q			<=			16'h0107;
		end
		32'h00007FF0: begin
				q			<=			16'h9793;
		end
		32'h00007FF2: begin
				q			<=			16'h0107;
		end
		32'h00007FF4: begin
				q			<=			16'hE7B3;
		end
		32'h00007FF6: begin
				q			<=			16'h01D7;
		end
		32'h00007FF8: begin
				q			<=			16'h2E23;
		end
		32'h00007FFA: begin
				q			<=			16'hFEFF;
		end
		32'h00007FFC: begin
				q			<=			16'hE8E3;
		end
		32'h00007FFE: begin
				q			<=			16'hFB12;
		end
		32'h00008000: begin
				q			<=			16'h2023;
		end
		32'h00008002: begin
				q			<=			16'h009F;
		end
		32'h00008004: begin
				q			<=			16'h5283;
		end
		32'h00008006: begin
				q			<=			16'h0026;
		end
		32'h00008008: begin
				q			<=			16'h8663;
		end
		32'h0000800A: begin
				q			<=			16'h0602;
		end
		32'h0000800C: begin
				q			<=			16'h2783;
		end
		32'h0000800E: begin
				q			<=			16'h0008;
		end
		32'h00008010: begin
				q			<=			16'h0E93;
		end
		32'h00008012: begin
				q			<=			16'h0008;
		end
		32'h00008014: begin
				q			<=			16'h8F13;
		end
		32'h00008016: begin
				q			<=			16'h0005;
		end
		32'h00008018: begin
				q			<=			16'h0F93;
		end
		32'h0000801A: begin
				q			<=			16'h0000;
		end
		32'h0000801C: begin
				q			<=			16'h2703;
		end
		32'h0000801E: begin
				q			<=			16'h000F;
		end
		32'h00008020: begin
				q			<=			16'hD383;
		end
		32'h00008022: begin
				q			<=			16'h002E;
		end
		32'h00008024: begin
				q			<=			16'hF7B3;
		end
		32'h00008026: begin
				q			<=			16'h00D7;
		end
		32'h00008028: begin
				q			<=			16'h7733;
		end
		32'h0000802A: begin
				q			<=			16'h00D7;
		end
		32'h0000802C: begin
				q			<=			16'h0733;
		end
		32'h0000802E: begin
				q			<=			16'h0257;
		end
		32'h00008030: begin
				q			<=			16'h8E93;
		end
		32'h00008032: begin
				q			<=			16'h004E;
		end
		32'h00008034: begin
				q			<=			16'h0F13;
		end
		32'h00008036: begin
				q			<=			16'h004F;
		end
		32'h00008038: begin
				q			<=			16'h0733;
		end
		32'h0000803A: begin
				q			<=			16'h0077;
		end
		32'h0000803C: begin
				q			<=			16'h0733;
		end
		32'h0000803E: begin
				q			<=			16'h01F7;
		end
		32'h00008040: begin
				q			<=			16'h1F93;
		end
		32'h00008042: begin
				q			<=			16'h0107;
		end
		32'h00008044: begin
				q			<=			16'hE7B3;
		end
		32'h00008046: begin
				q			<=			16'h00FF;
		end
		32'h00008048: begin
				q			<=			16'hAE23;
		end
		32'h0000804A: begin
				q			<=			16'hFEFE;
		end
		32'h0000804C: begin
				q			<=			16'h5783;
		end
		32'h0000804E: begin
				q			<=			16'hFFEF;
		end
		32'h00008050: begin
				q			<=			16'hAF83;
		end
		32'h00008052: begin
				q			<=			16'h000E;
		end
		32'h00008054: begin
				q			<=			16'h5713;
		end
		32'h00008056: begin
				q			<=			16'h0107;
		end
		32'h00008058: begin
				q			<=			16'h87B3;
		end
		32'h0000805A: begin
				q			<=			16'h0257;
		end
		32'h0000805C: begin
				q			<=			16'hFFB3;
		end
		32'h0000805E: begin
				q			<=			16'h00DF;
		end
		32'h00008060: begin
				q			<=			16'h87B3;
		end
		32'h00008062: begin
				q			<=			16'h01F7;
		end
		32'h00008064: begin
				q			<=			16'h87B3;
		end
		32'h00008066: begin
				q			<=			16'h00E7;
		end
		32'h00008068: begin
				q			<=			16'hDF93;
		end
		32'h0000806A: begin
				q			<=			16'h0107;
		end
		32'h0000806C: begin
				q			<=			16'h68E3;
		end
		32'h0000806E: begin
				q			<=			16'hFB1F;
		end
		32'h00008070: begin
				q			<=			16'hA023;
		end
		32'h00008072: begin
				q			<=			16'h00FE;
		end
		32'h00008074: begin
				q			<=			16'h0613;
		end
		32'h00008076: begin
				q			<=			16'h0046;
		end
		32'h00008078: begin
				q			<=			16'h0813;
		end
		32'h0000807A: begin
				q			<=			16'h0048;
		end
		32'h0000807C: begin
				q			<=			16'hF06F;
		end
		32'h0000807E: begin
				q			<=			16'hED9F;
		end
		32'h00008080: begin
				q			<=			16'h0413;
		end
		32'h00008082: begin
				q			<=			16'hFFF4;
		end
		32'h00008084: begin
				q			<=			16'hF06F;
		end
		32'h00008086: begin
				q			<=			16'hED5F;
		end
		32'h00008088: begin
				q			<=			16'h0113;
		end
		32'h0000808A: begin
				q			<=			16'hFE01;
		end
		32'h0000808C: begin
				q			<=			16'h2A23;
		end
		32'h0000808E: begin
				q			<=			16'h0091;
		end
		32'h00008090: begin
				q			<=			16'h2823;
		end
		32'h00008092: begin
				q			<=			16'h0121;
		end
		32'h00008094: begin
				q			<=			16'h2623;
		end
		32'h00008096: begin
				q			<=			16'h0131;
		end
		32'h00008098: begin
				q			<=			16'h2E23;
		end
		32'h0000809A: begin
				q			<=			16'h0011;
		end
		32'h0000809C: begin
				q			<=			16'h2C23;
		end
		32'h0000809E: begin
				q			<=			16'h0081;
		end
		32'h000080A0: begin
				q			<=			16'h2423;
		end
		32'h000080A2: begin
				q			<=			16'h0141;
		end
		32'h000080A4: begin
				q			<=			16'h7793;
		end
		32'h000080A6: begin
				q			<=			16'h0036;
		end
		32'h000080A8: begin
				q			<=			16'h0913;
		end
		32'h000080AA: begin
				q			<=			16'h0005;
		end
		32'h000080AC: begin
				q			<=			16'h0493;
		end
		32'h000080AE: begin
				q			<=			16'h0006;
		end
		32'h000080B0: begin
				q			<=			16'h8993;
		end
		32'h000080B2: begin
				q			<=			16'h0005;
		end
		32'h000080B4: begin
				q			<=			16'h8463;
		end
		32'h000080B6: begin
				q			<=			16'h0207;
		end
		32'h000080B8: begin
				q			<=			16'h8793;
		end
		32'h000080BA: begin
				q			<=			16'hFFF7;
		end
		32'h000080BC: begin
				q			<=			16'h7717;
		end
		32'h000080BE: begin
				q			<=			16'h0000;
		end
		32'h000080C0: begin
				q			<=			16'h0713;
		end
		32'h000080C2: begin
				q			<=			16'h4447;
		end
		32'h000080C4: begin
				q			<=			16'h9793;
		end
		32'h000080C6: begin
				q			<=			16'h0027;
		end
		32'h000080C8: begin
				q			<=			16'h07B3;
		end
		32'h000080CA: begin
				q			<=			16'h00F7;
		end
		32'h000080CC: begin
				q			<=			16'hA603;
		end
		32'h000080CE: begin
				q			<=			16'h0007;
		end
		32'h000080D0: begin
				q			<=			16'h0693;
		end
		32'h000080D2: begin
				q			<=			16'h0000;
		end
		32'h000080D4: begin
				q			<=			16'hF0EF;
		end
		32'h000080D6: begin
				q			<=			16'hA85F;
		end
		32'h000080D8: begin
				q			<=			16'h0993;
		end
		32'h000080DA: begin
				q			<=			16'h0005;
		end
		32'h000080DC: begin
				q			<=			16'hD493;
		end
		32'h000080DE: begin
				q			<=			16'h4024;
		end
		32'h000080E0: begin
				q			<=			16'h8663;
		end
		32'h000080E2: begin
				q			<=			16'h0804;
		end
		32'h000080E4: begin
				q			<=			16'h2403;
		end
		32'h000080E6: begin
				q			<=			16'h0489;
		end
		32'h000080E8: begin
				q			<=			16'h1E63;
		end
		32'h000080EA: begin
				q			<=			16'h0004;
		end
		32'h000080EC: begin
				q			<=			16'h0593;
		end
		32'h000080EE: begin
				q			<=			16'h2710;
		end
		32'h000080F0: begin
				q			<=			16'h0513;
		end
		32'h000080F2: begin
				q			<=			16'h0009;
		end
		32'h000080F4: begin
				q			<=			16'hF0EF;
		end
		32'h000080F6: begin
				q			<=			16'hD9DF;
		end
		32'h000080F8: begin
				q			<=			16'h2423;
		end
		32'h000080FA: begin
				q			<=			16'h04A9;
		end
		32'h000080FC: begin
				q			<=			16'h0413;
		end
		32'h000080FE: begin
				q			<=			16'h0005;
		end
		32'h00008100: begin
				q			<=			16'h2023;
		end
		32'h00008102: begin
				q			<=			16'h0005;
		end
		32'h00008104: begin
				q			<=			16'hF793;
		end
		32'h00008106: begin
				q			<=			16'h0014;
		end
		32'h00008108: begin
				q			<=			16'h8863;
		end
		32'h0000810A: begin
				q			<=			16'h0207;
		end
		32'h0000810C: begin
				q			<=			16'h8593;
		end
		32'h0000810E: begin
				q			<=			16'h0009;
		end
		32'h00008110: begin
				q			<=			16'h0613;
		end
		32'h00008112: begin
				q			<=			16'h0004;
		end
		32'h00008114: begin
				q			<=			16'h0513;
		end
		32'h00008116: begin
				q			<=			16'h0009;
		end
		32'h00008118: begin
				q			<=			16'h0097;
		end
		32'h0000811A: begin
				q			<=			16'h0000;
		end
		32'h0000811C: begin
				q			<=			16'h80E7;
		end
		32'h0000811E: begin
				q			<=			16'hDAC0;
		end
		32'h00008120: begin
				q			<=			16'h0A13;
		end
		32'h00008122: begin
				q			<=			16'h0005;
		end
		32'h00008124: begin
				q			<=			16'h8593;
		end
		32'h00008126: begin
				q			<=			16'h0009;
		end
		32'h00008128: begin
				q			<=			16'h0513;
		end
		32'h0000812A: begin
				q			<=			16'h0009;
		end
		32'h0000812C: begin
				q			<=			16'h0097;
		end
		32'h0000812E: begin
				q			<=			16'h0000;
		end
		32'h00008130: begin
				q			<=			16'h80E7;
		end
		32'h00008132: begin
				q			<=			16'hA080;
		end
		32'h00008134: begin
				q			<=			16'h0993;
		end
		32'h00008136: begin
				q			<=			16'h000A;
		end
		32'h00008138: begin
				q			<=			16'hD493;
		end
		32'h0000813A: begin
				q			<=			16'h4014;
		end
		32'h0000813C: begin
				q			<=			16'h8863;
		end
		32'h0000813E: begin
				q			<=			16'h0204;
		end
		32'h00008140: begin
				q			<=			16'h2503;
		end
		32'h00008142: begin
				q			<=			16'h0004;
		end
		32'h00008144: begin
				q			<=			16'h1063;
		end
		32'h00008146: begin
				q			<=			16'h0205;
		end
		32'h00008148: begin
				q			<=			16'h0613;
		end
		32'h0000814A: begin
				q			<=			16'h0004;
		end
		32'h0000814C: begin
				q			<=			16'h0593;
		end
		32'h0000814E: begin
				q			<=			16'h0004;
		end
		32'h00008150: begin
				q			<=			16'h0513;
		end
		32'h00008152: begin
				q			<=			16'h0009;
		end
		32'h00008154: begin
				q			<=			16'h0097;
		end
		32'h00008156: begin
				q			<=			16'h0000;
		end
		32'h00008158: begin
				q			<=			16'h80E7;
		end
		32'h0000815A: begin
				q			<=			16'hD700;
		end
		32'h0000815C: begin
				q			<=			16'h2023;
		end
		32'h0000815E: begin
				q			<=			16'h00A4;
		end
		32'h00008160: begin
				q			<=			16'h2023;
		end
		32'h00008162: begin
				q			<=			16'h0005;
		end
		32'h00008164: begin
				q			<=			16'h0413;
		end
		32'h00008166: begin
				q			<=			16'h0005;
		end
		32'h00008168: begin
				q			<=			16'hF06F;
		end
		32'h0000816A: begin
				q			<=			16'hF9DF;
		end
		32'h0000816C: begin
				q			<=			16'h2083;
		end
		32'h0000816E: begin
				q			<=			16'h01C1;
		end
		32'h00008170: begin
				q			<=			16'h2403;
		end
		32'h00008172: begin
				q			<=			16'h0181;
		end
		32'h00008174: begin
				q			<=			16'h8513;
		end
		32'h00008176: begin
				q			<=			16'h0009;
		end
		32'h00008178: begin
				q			<=			16'h2483;
		end
		32'h0000817A: begin
				q			<=			16'h0141;
		end
		32'h0000817C: begin
				q			<=			16'h2903;
		end
		32'h0000817E: begin
				q			<=			16'h0101;
		end
		32'h00008180: begin
				q			<=			16'h2983;
		end
		32'h00008182: begin
				q			<=			16'h00C1;
		end
		32'h00008184: begin
				q			<=			16'h2A03;
		end
		32'h00008186: begin
				q			<=			16'h0081;
		end
		32'h00008188: begin
				q			<=			16'h0113;
		end
		32'h0000818A: begin
				q			<=			16'h0201;
		end
		32'h0000818C: begin
				q			<=			16'h8067;
		end
		32'h0000818E: begin
				q			<=			16'h0000;
		end
		32'h00008190: begin
				q			<=			16'h0113;
		end
		32'h00008192: begin
				q			<=			16'hFD01;
		end
		32'h00008194: begin
				q			<=			16'h2223;
		end
		32'h00008196: begin
				q			<=			16'h0291;
		end
		32'h00008198: begin
				q			<=			16'h8493;
		end
		32'h0000819A: begin
				q			<=			16'h0005;
		end
		32'h0000819C: begin
				q			<=			16'h2E23;
		end
		32'h0000819E: begin
				q			<=			16'h0131;
		end
		32'h000081A0: begin
				q			<=			16'hA983;
		end
		32'h000081A2: begin
				q			<=			16'h0104;
		end
		32'h000081A4: begin
				q			<=			16'h2423;
		end
		32'h000081A6: begin
				q			<=			16'h0281;
		end
		32'h000081A8: begin
				q			<=			16'hA583;
		end
		32'h000081AA: begin
				q			<=			16'h0045;
		end
		32'h000081AC: begin
				q			<=			16'h5413;
		end
		32'h000081AE: begin
				q			<=			16'h4056;
		end
		32'h000081B0: begin
				q			<=			16'hA783;
		end
		32'h000081B2: begin
				q			<=			16'h0084;
		end
		32'h000081B4: begin
				q			<=			16'h09B3;
		end
		32'h000081B6: begin
				q			<=			16'h0134;
		end
		32'h000081B8: begin
				q			<=			16'h2023;
		end
		32'h000081BA: begin
				q			<=			16'h0321;
		end
		32'h000081BC: begin
				q			<=			16'h2A23;
		end
		32'h000081BE: begin
				q			<=			16'h0151;
		end
		32'h000081C0: begin
				q			<=			16'h2623;
		end
		32'h000081C2: begin
				q			<=			16'h0211;
		end
		32'h000081C4: begin
				q			<=			16'h2C23;
		end
		32'h000081C6: begin
				q			<=			16'h0141;
		end
		32'h000081C8: begin
				q			<=			16'h0A93;
		end
		32'h000081CA: begin
				q			<=			16'h0005;
		end
		32'h000081CC: begin
				q			<=			16'h8913;
		end
		32'h000081CE: begin
				q			<=			16'h0019;
		end
		32'h000081D0: begin
				q			<=			16'hC863;
		end
		32'h000081D2: begin
				q			<=			16'h0D27;
		end
		32'h000081D4: begin
				q			<=			16'h8513;
		end
		32'h000081D6: begin
				q			<=			16'h000A;
		end
		32'h000081D8: begin
				q			<=			16'h2623;
		end
		32'h000081DA: begin
				q			<=			16'h00C1;
		end
		32'h000081DC: begin
				q			<=			16'h0097;
		end
		32'h000081DE: begin
				q			<=			16'h0000;
		end
		32'h000081E0: begin
				q			<=			16'h80E7;
		end
		32'h000081E2: begin
				q			<=			16'h8B00;
		end
		32'h000081E4: begin
				q			<=			16'h2603;
		end
		32'h000081E6: begin
				q			<=			16'h00C1;
		end
		32'h000081E8: begin
				q			<=			16'h0793;
		end
		32'h000081EA: begin
				q			<=			16'h0145;
		end
		32'h000081EC: begin
				q			<=			16'h0A13;
		end
		32'h000081EE: begin
				q			<=			16'h0005;
		end
		32'h000081F0: begin
				q			<=			16'h8693;
		end
		32'h000081F2: begin
				q			<=			16'h0007;
		end
		32'h000081F4: begin
				q			<=			16'h0713;
		end
		32'h000081F6: begin
				q			<=			16'h0000;
		end
		32'h000081F8: begin
				q			<=			16'h8693;
		end
		32'h000081FA: begin
				q			<=			16'h0046;
		end
		32'h000081FC: begin
				q			<=			16'h4863;
		end
		32'h000081FE: begin
				q			<=			16'h0A87;
		end
		32'h00008200: begin
				q			<=			16'h5463;
		end
		32'h00008202: begin
				q			<=			16'h0004;
		end
		32'h00008204: begin
				q			<=			16'h0413;
		end
		32'h00008206: begin
				q			<=			16'h0000;
		end
		32'h00008208: begin
				q			<=			16'hA683;
		end
		32'h0000820A: begin
				q			<=			16'h0104;
		end
		32'h0000820C: begin
				q			<=			16'h1413;
		end
		32'h0000820E: begin
				q			<=			16'h0024;
		end
		32'h00008210: begin
				q			<=			16'h8733;
		end
		32'h00008212: begin
				q			<=			16'h0087;
		end
		32'h00008214: begin
				q			<=			16'h9693;
		end
		32'h00008216: begin
				q			<=			16'h0026;
		end
		32'h00008218: begin
				q			<=			16'h8793;
		end
		32'h0000821A: begin
				q			<=			16'h0144;
		end
		32'h0000821C: begin
				q			<=			16'h7613;
		end
		32'h0000821E: begin
				q			<=			16'h01F6;
		end
		32'h00008220: begin
				q			<=			16'h86B3;
		end
		32'h00008222: begin
				q			<=			16'h00D7;
		end
		32'h00008224: begin
				q			<=			16'h0A63;
		end
		32'h00008226: begin
				q			<=			16'h0806;
		end
		32'h00008228: begin
				q			<=			16'h0813;
		end
		32'h0000822A: begin
				q			<=			16'h0200;
		end
		32'h0000822C: begin
				q			<=			16'h0833;
		end
		32'h0000822E: begin
				q			<=			16'h40C8;
		end
		32'h00008230: begin
				q			<=			16'h0593;
		end
		32'h00008232: begin
				q			<=			16'h0000;
		end
		32'h00008234: begin
				q			<=			16'hA503;
		end
		32'h00008236: begin
				q			<=			16'h0007;
		end
		32'h00008238: begin
				q			<=			16'h0713;
		end
		32'h0000823A: begin
				q			<=			16'h0047;
		end
		32'h0000823C: begin
				q			<=			16'h8793;
		end
		32'h0000823E: begin
				q			<=			16'h0047;
		end
		32'h00008240: begin
				q			<=			16'h1533;
		end
		32'h00008242: begin
				q			<=			16'h00C5;
		end
		32'h00008244: begin
				q			<=			16'h65B3;
		end
		32'h00008246: begin
				q			<=			16'h00B5;
		end
		32'h00008248: begin
				q			<=			16'h2E23;
		end
		32'h0000824A: begin
				q			<=			16'hFEB7;
		end
		32'h0000824C: begin
				q			<=			16'hA583;
		end
		32'h0000824E: begin
				q			<=			16'hFFC7;
		end
		32'h00008250: begin
				q			<=			16'hD5B3;
		end
		32'h00008252: begin
				q			<=			16'h0105;
		end
		32'h00008254: begin
				q			<=			16'hE0E3;
		end
		32'h00008256: begin
				q			<=			16'hFED7;
		end
		32'h00008258: begin
				q			<=			16'h2023;
		end
		32'h0000825A: begin
				q			<=			16'h00B7;
		end
		32'h0000825C: begin
				q			<=			16'h8463;
		end
		32'h0000825E: begin
				q			<=			16'h0005;
		end
		32'h00008260: begin
				q			<=			16'h8913;
		end
		32'h00008262: begin
				q			<=			16'h0029;
		end
		32'h00008264: begin
				q			<=			16'h0913;
		end
		32'h00008266: begin
				q			<=			16'hFFF9;
		end
		32'h00008268: begin
				q			<=			16'h2823;
		end
		32'h0000826A: begin
				q			<=			16'h012A;
		end
		32'h0000826C: begin
				q			<=			16'h8513;
		end
		32'h0000826E: begin
				q			<=			16'h000A;
		end
		32'h00008270: begin
				q			<=			16'h8593;
		end
		32'h00008272: begin
				q			<=			16'h0004;
		end
		32'h00008274: begin
				q			<=			16'hF0EF;
		end
		32'h00008276: begin
				q			<=			16'h8C1F;
		end
		32'h00008278: begin
				q			<=			16'h2083;
		end
		32'h0000827A: begin
				q			<=			16'h02C1;
		end
		32'h0000827C: begin
				q			<=			16'h2403;
		end
		32'h0000827E: begin
				q			<=			16'h0281;
		end
		32'h00008280: begin
				q			<=			16'h0513;
		end
		32'h00008282: begin
				q			<=			16'h000A;
		end
		32'h00008284: begin
				q			<=			16'h2483;
		end
		32'h00008286: begin
				q			<=			16'h0241;
		end
		32'h00008288: begin
				q			<=			16'h2903;
		end
		32'h0000828A: begin
				q			<=			16'h0201;
		end
		32'h0000828C: begin
				q			<=			16'h2983;
		end
		32'h0000828E: begin
				q			<=			16'h01C1;
		end
		32'h00008290: begin
				q			<=			16'h2A03;
		end
		32'h00008292: begin
				q			<=			16'h0181;
		end
		32'h00008294: begin
				q			<=			16'h2A83;
		end
		32'h00008296: begin
				q			<=			16'h0141;
		end
		32'h00008298: begin
				q			<=			16'h0113;
		end
		32'h0000829A: begin
				q			<=			16'h0301;
		end
		32'h0000829C: begin
				q			<=			16'h8067;
		end
		32'h0000829E: begin
				q			<=			16'h0000;
		end
		32'h000082A0: begin
				q			<=			16'h8593;
		end
		32'h000082A2: begin
				q			<=			16'h0015;
		end
		32'h000082A4: begin
				q			<=			16'h9793;
		end
		32'h000082A6: begin
				q			<=			16'h0017;
		end
		32'h000082A8: begin
				q			<=			16'hF06F;
		end
		32'h000082AA: begin
				q			<=			16'hF29F;
		end
		32'h000082AC: begin
				q			<=			16'hAE23;
		end
		32'h000082AE: begin
				q			<=			16'hFE06;
		end
		32'h000082B0: begin
				q			<=			16'h0713;
		end
		32'h000082B2: begin
				q			<=			16'h0017;
		end
		32'h000082B4: begin
				q			<=			16'hF06F;
		end
		32'h000082B6: begin
				q			<=			16'hF45F;
		end
		32'h000082B8: begin
				q			<=			16'h8793;
		end
		32'h000082BA: begin
				q			<=			16'h0047;
		end
		32'h000082BC: begin
				q			<=			16'hA603;
		end
		32'h000082BE: begin
				q			<=			16'hFFC7;
		end
		32'h000082C0: begin
				q			<=			16'h0713;
		end
		32'h000082C2: begin
				q			<=			16'h0047;
		end
		32'h000082C4: begin
				q			<=			16'h2E23;
		end
		32'h000082C6: begin
				q			<=			16'hFEC7;
		end
		32'h000082C8: begin
				q			<=			16'hE8E3;
		end
		32'h000082CA: begin
				q			<=			16'hFED7;
		end
		32'h000082CC: begin
				q			<=			16'hF06F;
		end
		32'h000082CE: begin
				q			<=			16'hF99F;
		end
		32'h000082D0: begin
				q			<=			16'h2783;
		end
		32'h000082D2: begin
				q			<=			16'h0105;
		end
		32'h000082D4: begin
				q			<=			16'hA703;
		end
		32'h000082D6: begin
				q			<=			16'h0105;
		end
		32'h000082D8: begin
				q			<=			16'h87B3;
		end
		32'h000082DA: begin
				q			<=			16'h40E7;
		end
		32'h000082DC: begin
				q			<=			16'h9C63;
		end
		32'h000082DE: begin
				q			<=			16'h0207;
		end
		32'h000082E0: begin
				q			<=			16'h1713;
		end
		32'h000082E2: begin
				q			<=			16'h0027;
		end
		32'h000082E4: begin
				q			<=			16'h0513;
		end
		32'h000082E6: begin
				q			<=			16'h0145;
		end
		32'h000082E8: begin
				q			<=			16'h8593;
		end
		32'h000082EA: begin
				q			<=			16'h0145;
		end
		32'h000082EC: begin
				q			<=			16'h06B3;
		end
		32'h000082EE: begin
				q			<=			16'h00E5;
		end
		32'h000082F0: begin
				q			<=			16'h85B3;
		end
		32'h000082F2: begin
				q			<=			16'h00E5;
		end
		32'h000082F4: begin
				q			<=			16'h8693;
		end
		32'h000082F6: begin
				q			<=			16'hFFC6;
		end
		32'h000082F8: begin
				q			<=			16'h8593;
		end
		32'h000082FA: begin
				q			<=			16'hFFC5;
		end
		32'h000082FC: begin
				q			<=			16'hA603;
		end
		32'h000082FE: begin
				q			<=			16'h0006;
		end
		32'h00008300: begin
				q			<=			16'hA703;
		end
		32'h00008302: begin
				q			<=			16'h0005;
		end
		32'h00008304: begin
				q			<=			16'h0C63;
		end
		32'h00008306: begin
				q			<=			16'h00E6;
		end
		32'h00008308: begin
				q			<=			16'h0793;
		end
		32'h0000830A: begin
				q			<=			16'hFFF0;
		end
		32'h0000830C: begin
				q			<=			16'h6463;
		end
		32'h0000830E: begin
				q			<=			16'h00E6;
		end
		32'h00008310: begin
				q			<=			16'h0793;
		end
		32'h00008312: begin
				q			<=			16'h0010;
		end
		32'h00008314: begin
				q			<=			16'h8513;
		end
		32'h00008316: begin
				q			<=			16'h0007;
		end
		32'h00008318: begin
				q			<=			16'h8067;
		end
		32'h0000831A: begin
				q			<=			16'h0000;
		end
		32'h0000831C: begin
				q			<=			16'h6CE3;
		end
		32'h0000831E: begin
				q			<=			16'hFCD5;
		end
		32'h00008320: begin
				q			<=			16'hF06F;
		end
		32'h00008322: begin
				q			<=			16'hFF5F;
		end
		32'h00008324: begin
				q			<=			16'h0113;
		end
		32'h00008326: begin
				q			<=			16'hFE01;
		end
		32'h00008328: begin
				q			<=			16'h2A23;
		end
		32'h0000832A: begin
				q			<=			16'h0091;
		end
		32'h0000832C: begin
				q			<=			16'h8493;
		end
		32'h0000832E: begin
				q			<=			16'h0005;
		end
		32'h00008330: begin
				q			<=			16'h2623;
		end
		32'h00008332: begin
				q			<=			16'h0131;
		end
		32'h00008334: begin
				q			<=			16'h0593;
		end
		32'h00008336: begin
				q			<=			16'h0006;
		end
		32'h00008338: begin
				q			<=			16'h0993;
		end
		32'h0000833A: begin
				q			<=			16'h0005;
		end
		32'h0000833C: begin
				q			<=			16'h8513;
		end
		32'h0000833E: begin
				q			<=			16'h0004;
		end
		32'h00008340: begin
				q			<=			16'h2C23;
		end
		32'h00008342: begin
				q			<=			16'h0081;
		end
		32'h00008344: begin
				q			<=			16'h2E23;
		end
		32'h00008346: begin
				q			<=			16'h0011;
		end
		32'h00008348: begin
				q			<=			16'h2823;
		end
		32'h0000834A: begin
				q			<=			16'h0121;
		end
		32'h0000834C: begin
				q			<=			16'h0413;
		end
		32'h0000834E: begin
				q			<=			16'h0006;
		end
		32'h00008350: begin
				q			<=			16'h0097;
		end
		32'h00008352: begin
				q			<=			16'h0000;
		end
		32'h00008354: begin
				q			<=			16'h80E7;
		end
		32'h00008356: begin
				q			<=			16'hF800;
		end
		32'h00008358: begin
				q			<=			16'h1E63;
		end
		32'h0000835A: begin
				q			<=			16'h0205;
		end
		32'h0000835C: begin
				q			<=			16'h0593;
		end
		32'h0000835E: begin
				q			<=			16'h0000;
		end
		32'h00008360: begin
				q			<=			16'h8513;
		end
		32'h00008362: begin
				q			<=			16'h0009;
		end
		32'h00008364: begin
				q			<=			16'hF097;
		end
		32'h00008366: begin
				q			<=			16'hFFFF;
		end
		32'h00008368: begin
				q			<=			16'h80E7;
		end
		32'h0000836A: begin
				q			<=			16'h7280;
		end
		32'h0000836C: begin
				q			<=			16'h0793;
		end
		32'h0000836E: begin
				q			<=			16'h0010;
		end
		32'h00008370: begin
				q			<=			16'h2823;
		end
		32'h00008372: begin
				q			<=			16'h00F5;
		end
		32'h00008374: begin
				q			<=			16'h2A23;
		end
		32'h00008376: begin
				q			<=			16'h0005;
		end
		32'h00008378: begin
				q			<=			16'h2083;
		end
		32'h0000837A: begin
				q			<=			16'h01C1;
		end
		32'h0000837C: begin
				q			<=			16'h2403;
		end
		32'h0000837E: begin
				q			<=			16'h0181;
		end
		32'h00008380: begin
				q			<=			16'h2483;
		end
		32'h00008382: begin
				q			<=			16'h0141;
		end
		32'h00008384: begin
				q			<=			16'h2903;
		end
		32'h00008386: begin
				q			<=			16'h0101;
		end
		32'h00008388: begin
				q			<=			16'h2983;
		end
		32'h0000838A: begin
				q			<=			16'h00C1;
		end
		32'h0000838C: begin
				q			<=			16'h0113;
		end
		32'h0000838E: begin
				q			<=			16'h0201;
		end
		32'h00008390: begin
				q			<=			16'h8067;
		end
		32'h00008392: begin
				q			<=			16'h0000;
		end
		32'h00008394: begin
				q			<=			16'h0913;
		end
		32'h00008396: begin
				q			<=			16'h0010;
		end
		32'h00008398: begin
				q			<=			16'h4A63;
		end
		32'h0000839A: begin
				q			<=			16'h0005;
		end
		32'h0000839C: begin
				q			<=			16'h0793;
		end
		32'h0000839E: begin
				q			<=			16'h0004;
		end
		32'h000083A0: begin
				q			<=			16'h0913;
		end
		32'h000083A2: begin
				q			<=			16'h0000;
		end
		32'h000083A4: begin
				q			<=			16'h8413;
		end
		32'h000083A6: begin
				q			<=			16'h0004;
		end
		32'h000083A8: begin
				q			<=			16'h8493;
		end
		32'h000083AA: begin
				q			<=			16'h0007;
		end
		32'h000083AC: begin
				q			<=			16'h2583;
		end
		32'h000083AE: begin
				q			<=			16'h0044;
		end
		32'h000083B0: begin
				q			<=			16'h8513;
		end
		32'h000083B2: begin
				q			<=			16'h0009;
		end
		32'h000083B4: begin
				q			<=			16'hF097;
		end
		32'h000083B6: begin
				q			<=			16'hFFFF;
		end
		32'h000083B8: begin
				q			<=			16'h80E7;
		end
		32'h000083BA: begin
				q			<=			16'h6D80;
		end
		32'h000083BC: begin
				q			<=			16'h2303;
		end
		32'h000083BE: begin
				q			<=			16'h0104;
		end
		32'h000083C0: begin
				q			<=			16'hA883;
		end
		32'h000083C2: begin
				q			<=			16'h0104;
		end
		32'h000083C4: begin
				q			<=			16'h0613;
		end
		32'h000083C6: begin
				q			<=			16'h0144;
		end
		32'h000083C8: begin
				q			<=			16'h1E13;
		end
		32'h000083CA: begin
				q			<=			16'h0023;
		end
		32'h000083CC: begin
				q			<=			16'h8813;
		end
		32'h000083CE: begin
				q			<=			16'h0144;
		end
		32'h000083D0: begin
				q			<=			16'h9893;
		end
		32'h000083D2: begin
				q			<=			16'h0028;
		end
		32'h000083D4: begin
				q			<=			16'h0EB7;
		end
		32'h000083D6: begin
				q			<=			16'h0001;
		end
		32'h000083D8: begin
				q			<=			16'h2623;
		end
		32'h000083DA: begin
				q			<=			16'h0125;
		end
		32'h000083DC: begin
				q			<=			16'h0E33;
		end
		32'h000083DE: begin
				q			<=			16'h01C6;
		end
		32'h000083E0: begin
				q			<=			16'h08B3;
		end
		32'h000083E2: begin
				q			<=			16'h0118;
		end
		32'h000083E4: begin
				q			<=			16'h0693;
		end
		32'h000083E6: begin
				q			<=			16'h0145;
		end
		32'h000083E8: begin
				q			<=			16'h0F13;
		end
		32'h000083EA: begin
				q			<=			16'h0000;
		end
		32'h000083EC: begin
				q			<=			16'h8E93;
		end
		32'h000083EE: begin
				q			<=			16'hFFFE;
		end
		32'h000083F0: begin
				q			<=			16'h2703;
		end
		32'h000083F2: begin
				q			<=			16'h0006;
		end
		32'h000083F4: begin
				q			<=			16'h2F83;
		end
		32'h000083F6: begin
				q			<=			16'h0008;
		end
		32'h000083F8: begin
				q			<=			16'h8693;
		end
		32'h000083FA: begin
				q			<=			16'h0046;
		end
		32'h000083FC: begin
				q			<=			16'h75B3;
		end
		32'h000083FE: begin
				q			<=			16'h01D7;
		end
		32'h00008400: begin
				q			<=			16'hF7B3;
		end
		32'h00008402: begin
				q			<=			16'h01DF;
		end
		32'h00008404: begin
				q			<=			16'h85B3;
		end
		32'h00008406: begin
				q			<=			16'h01E5;
		end
		32'h00008408: begin
				q			<=			16'h85B3;
		end
		32'h0000840A: begin
				q			<=			16'h40F5;
		end
		32'h0000840C: begin
				q			<=			16'hDF93;
		end
		32'h0000840E: begin
				q			<=			16'h010F;
		end
		32'h00008410: begin
				q			<=			16'h5793;
		end
		32'h00008412: begin
				q			<=			16'h0107;
		end
		32'h00008414: begin
				q			<=			16'h87B3;
		end
		32'h00008416: begin
				q			<=			16'h41F7;
		end
		32'h00008418: begin
				q			<=			16'hD713;
		end
		32'h0000841A: begin
				q			<=			16'h4105;
		end
		32'h0000841C: begin
				q			<=			16'h87B3;
		end
		32'h0000841E: begin
				q			<=			16'h00E7;
		end
		32'h00008420: begin
				q			<=			16'hDF13;
		end
		32'h00008422: begin
				q			<=			16'h4107;
		end
		32'h00008424: begin
				q			<=			16'hF5B3;
		end
		32'h00008426: begin
				q			<=			16'h01D5;
		end
		32'h00008428: begin
				q			<=			16'h9793;
		end
		32'h0000842A: begin
				q			<=			16'h0107;
		end
		32'h0000842C: begin
				q			<=			16'hE7B3;
		end
		32'h0000842E: begin
				q			<=			16'h00B7;
		end
		32'h00008430: begin
				q			<=			16'h0813;
		end
		32'h00008432: begin
				q			<=			16'h0048;
		end
		32'h00008434: begin
				q			<=			16'hAE23;
		end
		32'h00008436: begin
				q			<=			16'hFEF6;
		end
		32'h00008438: begin
				q			<=			16'h0613;
		end
		32'h0000843A: begin
				q			<=			16'h0046;
		end
		32'h0000843C: begin
				q			<=			16'h6AE3;
		end
		32'h0000843E: begin
				q			<=			16'hFB18;
		end
		32'h00008440: begin
				q			<=			16'h05B7;
		end
		32'h00008442: begin
				q			<=			16'h0001;
		end
		32'h00008444: begin
				q			<=			16'h8593;
		end
		32'h00008446: begin
				q			<=			16'hFFF5;
		end
		32'h00008448: begin
				q			<=			16'h6C63;
		end
		32'h0000844A: begin
				q			<=			16'h01C6;
		end
		32'h0000844C: begin
				q			<=			16'h8693;
		end
		32'h0000844E: begin
				q			<=			16'hFFC6;
		end
		32'h00008450: begin
				q			<=			16'hA783;
		end
		32'h00008452: begin
				q			<=			16'h0006;
		end
		32'h00008454: begin
				q			<=			16'h8263;
		end
		32'h00008456: begin
				q			<=			16'h0407;
		end
		32'h00008458: begin
				q			<=			16'h2823;
		end
		32'h0000845A: begin
				q			<=			16'h0065;
		end
		32'h0000845C: begin
				q			<=			16'hF06F;
		end
		32'h0000845E: begin
				q			<=			16'hF1DF;
		end
		32'h00008460: begin
				q			<=			16'h2783;
		end
		32'h00008462: begin
				q			<=			16'h0006;
		end
		32'h00008464: begin
				q			<=			16'h8693;
		end
		32'h00008466: begin
				q			<=			16'h0046;
		end
		32'h00008468: begin
				q			<=			16'h0613;
		end
		32'h0000846A: begin
				q			<=			16'h0046;
		end
		32'h0000846C: begin
				q			<=			16'hF733;
		end
		32'h0000846E: begin
				q			<=			16'h00B7;
		end
		32'h00008470: begin
				q			<=			16'h0733;
		end
		32'h00008472: begin
				q			<=			16'h01E7;
		end
		32'h00008474: begin
				q			<=			16'h5813;
		end
		32'h00008476: begin
				q			<=			16'h4107;
		end
		32'h00008478: begin
				q			<=			16'hD793;
		end
		32'h0000847A: begin
				q			<=			16'h0107;
		end
		32'h0000847C: begin
				q			<=			16'h87B3;
		end
		32'h0000847E: begin
				q			<=			16'h0107;
		end
		32'h00008480: begin
				q			<=			16'hDF13;
		end
		32'h00008482: begin
				q			<=			16'h4107;
		end
		32'h00008484: begin
				q			<=			16'h7733;
		end
		32'h00008486: begin
				q			<=			16'h00B7;
		end
		32'h00008488: begin
				q			<=			16'h9793;
		end
		32'h0000848A: begin
				q			<=			16'h0107;
		end
		32'h0000848C: begin
				q			<=			16'hE7B3;
		end
		32'h0000848E: begin
				q			<=			16'h00E7;
		end
		32'h00008490: begin
				q			<=			16'hAE23;
		end
		32'h00008492: begin
				q			<=			16'hFEF6;
		end
		32'h00008494: begin
				q			<=			16'hF06F;
		end
		32'h00008496: begin
				q			<=			16'hFB5F;
		end
		32'h00008498: begin
				q			<=			16'h0313;
		end
		32'h0000849A: begin
				q			<=			16'hFFF3;
		end
		32'h0000849C: begin
				q			<=			16'hF06F;
		end
		32'h0000849E: begin
				q			<=			16'hFB1F;
		end
		32'h000084A0: begin
				q			<=			16'h07B7;
		end
		32'h000084A2: begin
				q			<=			16'h7FF0;
		end
		32'h000084A4: begin
				q			<=			16'hF5B3;
		end
		32'h000084A6: begin
				q			<=			16'h00B7;
		end
		32'h000084A8: begin
				q			<=			16'h07B7;
		end
		32'h000084AA: begin
				q			<=			16'hFCC0;
		end
		32'h000084AC: begin
				q			<=			16'h85B3;
		end
		32'h000084AE: begin
				q			<=			16'h00F5;
		end
		32'h000084B0: begin
				q			<=			16'h5863;
		end
		32'h000084B2: begin
				q			<=			16'h00B0;
		end
		32'h000084B4: begin
				q			<=			16'h0793;
		end
		32'h000084B6: begin
				q			<=			16'h0000;
		end
		32'h000084B8: begin
				q			<=			16'h8513;
		end
		32'h000084BA: begin
				q			<=			16'h0007;
		end
		32'h000084BC: begin
				q			<=			16'h8067;
		end
		32'h000084BE: begin
				q			<=			16'h0000;
		end
		32'h000084C0: begin
				q			<=			16'h05B3;
		end
		32'h000084C2: begin
				q			<=			16'h40B0;
		end
		32'h000084C4: begin
				q			<=			16'hD793;
		end
		32'h000084C6: begin
				q			<=			16'h4145;
		end
		32'h000084C8: begin
				q			<=			16'h0713;
		end
		32'h000084CA: begin
				q			<=			16'h0130;
		end
		32'h000084CC: begin
				q			<=			16'h4863;
		end
		32'h000084CE: begin
				q			<=			16'h00F7;
		end
		32'h000084D0: begin
				q			<=			16'h05B7;
		end
		32'h000084D2: begin
				q			<=			16'h0008;
		end
		32'h000084D4: begin
				q			<=			16'hD5B3;
		end
		32'h000084D6: begin
				q			<=			16'h40F5;
		end
		32'h000084D8: begin
				q			<=			16'hF06F;
		end
		32'h000084DA: begin
				q			<=			16'hFDDF;
		end
		32'h000084DC: begin
				q			<=			16'h8793;
		end
		32'h000084DE: begin
				q			<=			16'hFEC7;
		end
		32'h000084E0: begin
				q			<=			16'h0693;
		end
		32'h000084E2: begin
				q			<=			16'h01E0;
		end
		32'h000084E4: begin
				q			<=			16'h0593;
		end
		32'h000084E6: begin
				q			<=			16'h0000;
		end
		32'h000084E8: begin
				q			<=			16'h0713;
		end
		32'h000084EA: begin
				q			<=			16'h0010;
		end
		32'h000084EC: begin
				q			<=			16'hC663;
		end
		32'h000084EE: begin
				q			<=			16'h00F6;
		end
		32'h000084F0: begin
				q			<=			16'hC793;
		end
		32'h000084F2: begin
				q			<=			16'hFFF7;
		end
		32'h000084F4: begin
				q			<=			16'h1733;
		end
		32'h000084F6: begin
				q			<=			16'h00F7;
		end
		32'h000084F8: begin
				q			<=			16'h0793;
		end
		32'h000084FA: begin
				q			<=			16'h0007;
		end
		32'h000084FC: begin
				q			<=			16'hF06F;
		end
		32'h000084FE: begin
				q			<=			16'hFBDF;
		end
		32'h00008500: begin
				q			<=			16'h0113;
		end
		32'h00008502: begin
				q			<=			16'hFD01;
		end
		32'h00008504: begin
				q			<=			16'h2223;
		end
		32'h00008506: begin
				q			<=			16'h0291;
		end
		32'h00008508: begin
				q			<=			16'h2483;
		end
		32'h0000850A: begin
				q			<=			16'h0105;
		end
		32'h0000850C: begin
				q			<=			16'h2E23;
		end
		32'h0000850E: begin
				q			<=			16'h0131;
		end
		32'h00008510: begin
				q			<=			16'h0993;
		end
		32'h00008512: begin
				q			<=			16'h0145;
		end
		32'h00008514: begin
				q			<=			16'h9493;
		end
		32'h00008516: begin
				q			<=			16'h0024;
		end
		32'h00008518: begin
				q			<=			16'h84B3;
		end
		32'h0000851A: begin
				q			<=			16'h0099;
		end
		32'h0000851C: begin
				q			<=			16'h2423;
		end
		32'h0000851E: begin
				q			<=			16'h0281;
		end
		32'h00008520: begin
				q			<=			16'hA403;
		end
		32'h00008522: begin
				q			<=			16'hFFC4;
		end
		32'h00008524: begin
				q			<=			16'h2023;
		end
		32'h00008526: begin
				q			<=			16'h0321;
		end
		32'h00008528: begin
				q			<=			16'h2623;
		end
		32'h0000852A: begin
				q			<=			16'h00B1;
		end
		32'h0000852C: begin
				q			<=			16'h0513;
		end
		32'h0000852E: begin
				q			<=			16'h0004;
		end
		32'h00008530: begin
				q			<=			16'h2623;
		end
		32'h00008532: begin
				q			<=			16'h0211;
		end
		32'h00008534: begin
				q			<=			16'h0097;
		end
		32'h00008536: begin
				q			<=			16'h0000;
		end
		32'h00008538: begin
				q			<=			16'h80E7;
		end
		32'h0000853A: begin
				q			<=			16'h8380;
		end
		32'h0000853C: begin
				q			<=			16'h2583;
		end
		32'h0000853E: begin
				q			<=			16'h00C1;
		end
		32'h00008540: begin
				q			<=			16'h0793;
		end
		32'h00008542: begin
				q			<=			16'h0200;
		end
		32'h00008544: begin
				q			<=			16'h87B3;
		end
		32'h00008546: begin
				q			<=			16'h40A7;
		end
		32'h00008548: begin
				q			<=			16'hA023;
		end
		32'h0000854A: begin
				q			<=			16'h00F5;
		end
		32'h0000854C: begin
				q			<=			16'h0793;
		end
		32'h0000854E: begin
				q			<=			16'h00A0;
		end
		32'h00008550: begin
				q			<=			16'h8913;
		end
		32'h00008552: begin
				q			<=			16'hFFC4;
		end
		32'h00008554: begin
				q			<=			16'hCC63;
		end
		32'h00008556: begin
				q			<=			16'h04A7;
		end
		32'h00008558: begin
				q			<=			16'h0793;
		end
		32'h0000855A: begin
				q			<=			16'h00B0;
		end
		32'h0000855C: begin
				q			<=			16'h87B3;
		end
		32'h0000855E: begin
				q			<=			16'h40A7;
		end
		32'h00008560: begin
				q			<=			16'h0737;
		end
		32'h00008562: begin
				q			<=			16'h3FF0;
		end
		32'h00008564: begin
				q			<=			16'h56B3;
		end
		32'h00008566: begin
				q			<=			16'h00F4;
		end
		32'h00008568: begin
				q			<=			16'hE6B3;
		end
		32'h0000856A: begin
				q			<=			16'h00E6;
		end
		32'h0000856C: begin
				q			<=			16'h0713;
		end
		32'h0000856E: begin
				q			<=			16'h0000;
		end
		32'h00008570: begin
				q			<=			16'hF463;
		end
		32'h00008572: begin
				q			<=			16'h0129;
		end
		32'h00008574: begin
				q			<=			16'hA703;
		end
		32'h00008576: begin
				q			<=			16'hFF84;
		end
		32'h00008578: begin
				q			<=			16'h0513;
		end
		32'h0000857A: begin
				q			<=			16'h0155;
		end
		32'h0000857C: begin
				q			<=			16'h1533;
		end
		32'h0000857E: begin
				q			<=			16'h00A4;
		end
		32'h00008580: begin
				q			<=			16'h57B3;
		end
		32'h00008582: begin
				q			<=			16'h00F7;
		end
		32'h00008584: begin
				q			<=			16'h67B3;
		end
		32'h00008586: begin
				q			<=			16'h00F5;
		end
		32'h00008588: begin
				q			<=			16'h2083;
		end
		32'h0000858A: begin
				q			<=			16'h02C1;
		end
		32'h0000858C: begin
				q			<=			16'h2403;
		end
		32'h0000858E: begin
				q			<=			16'h0281;
		end
		32'h00008590: begin
				q			<=			16'h2483;
		end
		32'h00008592: begin
				q			<=			16'h0241;
		end
		32'h00008594: begin
				q			<=			16'h2903;
		end
		32'h00008596: begin
				q			<=			16'h0201;
		end
		32'h00008598: begin
				q			<=			16'h2983;
		end
		32'h0000859A: begin
				q			<=			16'h01C1;
		end
		32'h0000859C: begin
				q			<=			16'h8513;
		end
		32'h0000859E: begin
				q			<=			16'h0007;
		end
		32'h000085A0: begin
				q			<=			16'h8593;
		end
		32'h000085A2: begin
				q			<=			16'h0006;
		end
		32'h000085A4: begin
				q			<=			16'h0113;
		end
		32'h000085A6: begin
				q			<=			16'h0301;
		end
		32'h000085A8: begin
				q			<=			16'h8067;
		end
		32'h000085AA: begin
				q			<=			16'h0000;
		end
		32'h000085AC: begin
				q			<=			16'h0793;
		end
		32'h000085AE: begin
				q			<=			16'h0000;
		end
		32'h000085B0: begin
				q			<=			16'hF663;
		end
		32'h000085B2: begin
				q			<=			16'h0129;
		end
		32'h000085B4: begin
				q			<=			16'hA783;
		end
		32'h000085B6: begin
				q			<=			16'hFF84;
		end
		32'h000085B8: begin
				q			<=			16'h8913;
		end
		32'h000085BA: begin
				q			<=			16'hFF84;
		end
		32'h000085BC: begin
				q			<=			16'h0513;
		end
		32'h000085BE: begin
				q			<=			16'hFF55;
		end
		32'h000085C0: begin
				q			<=			16'h0E63;
		end
		32'h000085C2: begin
				q			<=			16'h0205;
		end
		32'h000085C4: begin
				q			<=			16'h0713;
		end
		32'h000085C6: begin
				q			<=			16'h0200;
		end
		32'h000085C8: begin
				q			<=			16'h0633;
		end
		32'h000085CA: begin
				q			<=			16'h40A7;
		end
		32'h000085CC: begin
				q			<=			16'h1433;
		end
		32'h000085CE: begin
				q			<=			16'h00A4;
		end
		32'h000085D0: begin
				q			<=			16'h0737;
		end
		32'h000085D2: begin
				q			<=			16'h3FF0;
		end
		32'h000085D4: begin
				q			<=			16'h6433;
		end
		32'h000085D6: begin
				q			<=			16'h00E4;
		end
		32'h000085D8: begin
				q			<=			16'hD6B3;
		end
		32'h000085DA: begin
				q			<=			16'h00C7;
		end
		32'h000085DC: begin
				q			<=			16'h66B3;
		end
		32'h000085DE: begin
				q			<=			16'h00D4;
		end
		32'h000085E0: begin
				q			<=			16'h0713;
		end
		32'h000085E2: begin
				q			<=			16'h0000;
		end
		32'h000085E4: begin
				q			<=			16'hF463;
		end
		32'h000085E6: begin
				q			<=			16'h0129;
		end
		32'h000085E8: begin
				q			<=			16'h2703;
		end
		32'h000085EA: begin
				q			<=			16'hFFC9;
		end
		32'h000085EC: begin
				q			<=			16'h97B3;
		end
		32'h000085EE: begin
				q			<=			16'h00A7;
		end
		32'h000085F0: begin
				q			<=			16'h5733;
		end
		32'h000085F2: begin
				q			<=			16'h00C7;
		end
		32'h000085F4: begin
				q			<=			16'hE7B3;
		end
		32'h000085F6: begin
				q			<=			16'h00E7;
		end
		32'h000085F8: begin
				q			<=			16'hF06F;
		end
		32'h000085FA: begin
				q			<=			16'hF91F;
		end
		32'h000085FC: begin
				q			<=			16'h06B7;
		end
		32'h000085FE: begin
				q			<=			16'h3FF0;
		end
		32'h00008600: begin
				q			<=			16'h66B3;
		end
		32'h00008602: begin
				q			<=			16'h00D4;
		end
		32'h00008604: begin
				q			<=			16'hF06F;
		end
		32'h00008606: begin
				q			<=			16'hF85F;
		end
		32'h00008608: begin
				q			<=			16'h0113;
		end
		32'h0000860A: begin
				q			<=			16'hFD01;
		end
		32'h0000860C: begin
				q			<=			16'h2423;
		end
		32'h0000860E: begin
				q			<=			16'h0281;
		end
		32'h00008610: begin
				q			<=			16'h8413;
		end
		32'h00008612: begin
				q			<=			16'h0005;
		end
		32'h00008614: begin
				q			<=			16'h0593;
		end
		32'h00008616: begin
				q			<=			16'h0010;
		end
		32'h00008618: begin
				q			<=			16'h2223;
		end
		32'h0000861A: begin
				q			<=			16'h0291;
		end
		32'h0000861C: begin
				q			<=			16'h2023;
		end
		32'h0000861E: begin
				q			<=			16'h0321;
		end
		32'h00008620: begin
				q			<=			16'h0493;
		end
		32'h00008622: begin
				q			<=			16'h0006;
		end
		32'h00008624: begin
				q			<=			16'h2E23;
		end
		32'h00008626: begin
				q			<=			16'h0131;
		end
		32'h00008628: begin
				q			<=			16'h2C23;
		end
		32'h0000862A: begin
				q			<=			16'h0141;
		end
		32'h0000862C: begin
				q			<=			16'h0913;
		end
		32'h0000862E: begin
				q			<=			16'h0007;
		end
		32'h00008630: begin
				q			<=			16'h2623;
		end
		32'h00008632: begin
				q			<=			16'h0211;
		end
		32'h00008634: begin
				q			<=			16'h8A13;
		end
		32'h00008636: begin
				q			<=			16'h0006;
		end
		32'h00008638: begin
				q			<=			16'hF0EF;
		end
		32'h0000863A: begin
				q			<=			16'hC54F;
		end
		32'h0000863C: begin
				q			<=			16'h0737;
		end
		32'h0000863E: begin
				q			<=			16'h0010;
		end
		32'h00008640: begin
				q			<=			16'h0793;
		end
		32'h00008642: begin
				q			<=			16'hFFF7;
		end
		32'h00008644: begin
				q			<=			16'hF7B3;
		end
		32'h00008646: begin
				q			<=			16'h0097;
		end
		32'h00008648: begin
				q			<=			16'hD493;
		end
		32'h0000864A: begin
				q			<=			16'h0144;
		end
		32'h0000864C: begin
				q			<=			16'hF493;
		end
		32'h0000864E: begin
				q			<=			16'h7FF4;
		end
		32'h00008650: begin
				q			<=			16'h0993;
		end
		32'h00008652: begin
				q			<=			16'h0005;
		end
		32'h00008654: begin
				q			<=			16'h9C63;
		end
		32'h00008656: begin
				q			<=			16'h0804;
		end
		32'h00008658: begin
				q			<=			16'h2623;
		end
		32'h0000865A: begin
				q			<=			16'h00F1;
		end
		32'h0000865C: begin
				q			<=			16'h0063;
		end
		32'h0000865E: begin
				q			<=			16'h0A04;
		end
		32'h00008660: begin
				q			<=			16'h0513;
		end
		32'h00008662: begin
				q			<=			16'h0081;
		end
		32'h00008664: begin
				q			<=			16'h2423;
		end
		32'h00008666: begin
				q			<=			16'h0081;
		end
		32'h00008668: begin
				q			<=			16'hF097;
		end
		32'h0000866A: begin
				q			<=			16'hFFFF;
		end
		32'h0000866C: begin
				q			<=			16'h80E7;
		end
		32'h0000866E: begin
				q			<=			16'h7780;
		end
		32'h00008670: begin
				q			<=			16'h2683;
		end
		32'h00008672: begin
				q			<=			16'h0081;
		end
		32'h00008674: begin
				q			<=			16'h0063;
		end
		32'h00008676: begin
				q			<=			16'h0805;
		end
		32'h00008678: begin
				q			<=			16'h2703;
		end
		32'h0000867A: begin
				q			<=			16'h00C1;
		end
		32'h0000867C: begin
				q			<=			16'h0793;
		end
		32'h0000867E: begin
				q			<=			16'h0200;
		end
		32'h00008680: begin
				q			<=			16'h87B3;
		end
		32'h00008682: begin
				q			<=			16'h40A7;
		end
		32'h00008684: begin
				q			<=			16'h17B3;
		end
		32'h00008686: begin
				q			<=			16'h00F7;
		end
		32'h00008688: begin
				q			<=			16'hE7B3;
		end
		32'h0000868A: begin
				q			<=			16'h00D7;
		end
		32'h0000868C: begin
				q			<=			16'h5733;
		end
		32'h0000868E: begin
				q			<=			16'h00A7;
		end
		32'h00008690: begin
				q			<=			16'hAA23;
		end
		32'h00008692: begin
				q			<=			16'h00F9;
		end
		32'h00008694: begin
				q			<=			16'h2623;
		end
		32'h00008696: begin
				q			<=			16'h00E1;
		end
		32'h00008698: begin
				q			<=			16'h2403;
		end
		32'h0000869A: begin
				q			<=			16'h00C1;
		end
		32'h0000869C: begin
				q			<=			16'hAC23;
		end
		32'h0000869E: begin
				q			<=			16'h0089;
		end
		32'h000086A0: begin
				q			<=			16'h3433;
		end
		32'h000086A2: begin
				q			<=			16'h0080;
		end
		32'h000086A4: begin
				q			<=			16'h0413;
		end
		32'h000086A6: begin
				q			<=			16'h0014;
		end
		32'h000086A8: begin
				q			<=			16'hA823;
		end
		32'h000086AA: begin
				q			<=			16'h0089;
		end
		32'h000086AC: begin
				q			<=			16'h8C63;
		end
		32'h000086AE: begin
				q			<=			16'h0604;
		end
		32'h000086B0: begin
				q			<=			16'h8493;
		end
		32'h000086B2: begin
				q			<=			16'hBCD4;
		end
		32'h000086B4: begin
				q			<=			16'h84B3;
		end
		32'h000086B6: begin
				q			<=			16'h00A4;
		end
		32'h000086B8: begin
				q			<=			16'h0793;
		end
		32'h000086BA: begin
				q			<=			16'h0350;
		end
		32'h000086BC: begin
				q			<=			16'h2023;
		end
		32'h000086BE: begin
				q			<=			16'h009A;
		end
		32'h000086C0: begin
				q			<=			16'h8533;
		end
		32'h000086C2: begin
				q			<=			16'h40A7;
		end
		32'h000086C4: begin
				q			<=			16'h2023;
		end
		32'h000086C6: begin
				q			<=			16'h00A9;
		end
		32'h000086C8: begin
				q			<=			16'h2083;
		end
		32'h000086CA: begin
				q			<=			16'h02C1;
		end
		32'h000086CC: begin
				q			<=			16'h2403;
		end
		32'h000086CE: begin
				q			<=			16'h0281;
		end
		32'h000086D0: begin
				q			<=			16'h8513;
		end
		32'h000086D2: begin
				q			<=			16'h0009;
		end
		32'h000086D4: begin
				q			<=			16'h2483;
		end
		32'h000086D6: begin
				q			<=			16'h0241;
		end
		32'h000086D8: begin
				q			<=			16'h2903;
		end
		32'h000086DA: begin
				q			<=			16'h0201;
		end
		32'h000086DC: begin
				q			<=			16'h2983;
		end
		32'h000086DE: begin
				q			<=			16'h01C1;
		end
		32'h000086E0: begin
				q			<=			16'h2A03;
		end
		32'h000086E2: begin
				q			<=			16'h0181;
		end
		32'h000086E4: begin
				q			<=			16'h0113;
		end
		32'h000086E6: begin
				q			<=			16'h0301;
		end
		32'h000086E8: begin
				q			<=			16'h8067;
		end
		32'h000086EA: begin
				q			<=			16'h0000;
		end
		32'h000086EC: begin
				q			<=			16'hE7B3;
		end
		32'h000086EE: begin
				q			<=			16'h00E7;
		end
		32'h000086F0: begin
				q			<=			16'hF06F;
		end
		32'h000086F2: begin
				q			<=			16'hF69F;
		end
		32'h000086F4: begin
				q			<=			16'hAA23;
		end
		32'h000086F6: begin
				q			<=			16'h00D9;
		end
		32'h000086F8: begin
				q			<=			16'hF06F;
		end
		32'h000086FA: begin
				q			<=			16'hFA1F;
		end
		32'h000086FC: begin
				q			<=			16'h0513;
		end
		32'h000086FE: begin
				q			<=			16'h00C1;
		end
		32'h00008700: begin
				q			<=			16'hF097;
		end
		32'h00008702: begin
				q			<=			16'hFFFF;
		end
		32'h00008704: begin
				q			<=			16'h80E7;
		end
		32'h00008706: begin
				q			<=			16'h6E00;
		end
		32'h00008708: begin
				q			<=			16'h2783;
		end
		32'h0000870A: begin
				q			<=			16'h00C1;
		end
		32'h0000870C: begin
				q			<=			16'h0513;
		end
		32'h0000870E: begin
				q			<=			16'h0205;
		end
		32'h00008710: begin
				q			<=			16'h0413;
		end
		32'h00008712: begin
				q			<=			16'h0010;
		end
		32'h00008714: begin
				q			<=			16'hAA23;
		end
		32'h00008716: begin
				q			<=			16'h00F9;
		end
		32'h00008718: begin
				q			<=			16'h0793;
		end
		32'h0000871A: begin
				q			<=			16'h0010;
		end
		32'h0000871C: begin
				q			<=			16'hA823;
		end
		32'h0000871E: begin
				q			<=			16'h00F9;
		end
		32'h00008720: begin
				q			<=			16'hF06F;
		end
		32'h00008722: begin
				q			<=			16'hF8DF;
		end
		32'h00008724: begin
				q			<=			16'h1793;
		end
		32'h00008726: begin
				q			<=			16'h0024;
		end
		32'h00008728: begin
				q			<=			16'h0513;
		end
		32'h0000872A: begin
				q			<=			16'hBCE5;
		end
		32'h0000872C: begin
				q			<=			16'h87B3;
		end
		32'h0000872E: begin
				q			<=			16'h00F9;
		end
		32'h00008730: begin
				q			<=			16'h2023;
		end
		32'h00008732: begin
				q			<=			16'h00AA;
		end
		32'h00008734: begin
				q			<=			16'hA503;
		end
		32'h00008736: begin
				q			<=			16'h0107;
		end
		32'h00008738: begin
				q			<=			16'h1413;
		end
		32'h0000873A: begin
				q			<=			16'h0054;
		end
		32'h0000873C: begin
				q			<=			16'hF0EF;
		end
		32'h0000873E: begin
				q			<=			16'hE30F;
		end
		32'h00008740: begin
				q			<=			16'h0433;
		end
		32'h00008742: begin
				q			<=			16'h40A4;
		end
		32'h00008744: begin
				q			<=			16'h2023;
		end
		32'h00008746: begin
				q			<=			16'h0089;
		end
		32'h00008748: begin
				q			<=			16'hF06F;
		end
		32'h0000874A: begin
				q			<=			16'hF81F;
		end
		32'h0000874C: begin
				q			<=			16'h0113;
		end
		32'h0000874E: begin
				q			<=			16'hFD01;
		end
		32'h00008750: begin
				q			<=			16'h2023;
		end
		32'h00008752: begin
				q			<=			16'h0321;
		end
		32'h00008754: begin
				q			<=			16'h8913;
		end
		32'h00008756: begin
				q			<=			16'h0005;
		end
		32'h00008758: begin
				q			<=			16'h0593;
		end
		32'h0000875A: begin
				q			<=			16'h0081;
		end
		32'h0000875C: begin
				q			<=			16'h2623;
		end
		32'h0000875E: begin
				q			<=			16'h0211;
		end
		32'h00008760: begin
				q			<=			16'h2423;
		end
		32'h00008762: begin
				q			<=			16'h0281;
		end
		32'h00008764: begin
				q			<=			16'h2223;
		end
		32'h00008766: begin
				q			<=			16'h0291;
		end
		32'h00008768: begin
				q			<=			16'h2E23;
		end
		32'h0000876A: begin
				q			<=			16'h0131;
		end
		32'h0000876C: begin
				q			<=			16'h2C23;
		end
		32'h0000876E: begin
				q			<=			16'h0141;
		end
		32'h00008770: begin
				q			<=			16'h0A13;
		end
		32'h00008772: begin
				q			<=			16'h0005;
		end
		32'h00008774: begin
				q			<=			16'hF0EF;
		end
		32'h00008776: begin
				q			<=			16'hD8DF;
		end
		32'h00008778: begin
				q			<=			16'h0993;
		end
		32'h0000877A: begin
				q			<=			16'h0005;
		end
		32'h0000877C: begin
				q			<=			16'h8493;
		end
		32'h0000877E: begin
				q			<=			16'h0005;
		end
		32'h00008780: begin
				q			<=			16'h8413;
		end
		32'h00008782: begin
				q			<=			16'h0005;
		end
		32'h00008784: begin
				q			<=			16'h0513;
		end
		32'h00008786: begin
				q			<=			16'h0009;
		end
		32'h00008788: begin
				q			<=			16'h0593;
		end
		32'h0000878A: begin
				q			<=			16'h00C1;
		end
		32'h0000878C: begin
				q			<=			16'hF0EF;
		end
		32'h0000878E: begin
				q			<=			16'hD75F;
		end
		32'h00008790: begin
				q			<=			16'h2783;
		end
		32'h00008792: begin
				q			<=			16'h0109;
		end
		32'h00008794: begin
				q			<=			16'h2703;
		end
		32'h00008796: begin
				q			<=			16'h010A;
		end
		32'h00008798: begin
				q			<=			16'h2683;
		end
		32'h0000879A: begin
				q			<=			16'h0081;
		end
		32'h0000879C: begin
				q			<=			16'h0733;
		end
		32'h0000879E: begin
				q			<=			16'h40F7;
		end
		32'h000087A0: begin
				q			<=			16'h2783;
		end
		32'h000087A2: begin
				q			<=			16'h00C1;
		end
		32'h000087A4: begin
				q			<=			16'h1713;
		end
		32'h000087A6: begin
				q			<=			16'h0057;
		end
		32'h000087A8: begin
				q			<=			16'h86B3;
		end
		32'h000087AA: begin
				q			<=			16'h40F6;
		end
		32'h000087AC: begin
				q			<=			16'h07B3;
		end
		32'h000087AE: begin
				q			<=			16'h00D7;
		end
		32'h000087B0: begin
				q			<=			16'h5663;
		end
		32'h000087B2: begin
				q			<=			16'h04F0;
		end
		32'h000087B4: begin
				q			<=			16'h9793;
		end
		32'h000087B6: begin
				q			<=			16'h0147;
		end
		32'h000087B8: begin
				q			<=			16'h8613;
		end
		32'h000087BA: begin
				q			<=			16'h0005;
		end
		32'h000087BC: begin
				q			<=			16'h8433;
		end
		32'h000087BE: begin
				q			<=			16'h0097;
		end
		32'h000087C0: begin
				q			<=			16'h0713;
		end
		32'h000087C2: begin
				q			<=			16'h0006;
		end
		32'h000087C4: begin
				q			<=			16'h0593;
		end
		32'h000087C6: begin
				q			<=			16'h0004;
		end
		32'h000087C8: begin
				q			<=			16'h0613;
		end
		32'h000087CA: begin
				q			<=			16'h0005;
		end
		32'h000087CC: begin
				q			<=			16'h0693;
		end
		32'h000087CE: begin
				q			<=			16'h0007;
		end
		32'h000087D0: begin
				q			<=			16'h8513;
		end
		32'h000087D2: begin
				q			<=			16'h0009;
		end
		32'h000087D4: begin
				q			<=			16'h3097;
		end
		32'h000087D6: begin
				q			<=			16'h0000;
		end
		32'h000087D8: begin
				q			<=			16'h80E7;
		end
		32'h000087DA: begin
				q			<=			16'hB240;
		end
		32'h000087DC: begin
				q			<=			16'h2083;
		end
		32'h000087DE: begin
				q			<=			16'h02C1;
		end
		32'h000087E0: begin
				q			<=			16'h2403;
		end
		32'h000087E2: begin
				q			<=			16'h0281;
		end
		32'h000087E4: begin
				q			<=			16'h2483;
		end
		32'h000087E6: begin
				q			<=			16'h0241;
		end
		32'h000087E8: begin
				q			<=			16'h2903;
		end
		32'h000087EA: begin
				q			<=			16'h0201;
		end
		32'h000087EC: begin
				q			<=			16'h2983;
		end
		32'h000087EE: begin
				q			<=			16'h01C1;
		end
		32'h000087F0: begin
				q			<=			16'h2A03;
		end
		32'h000087F2: begin
				q			<=			16'h0181;
		end
		32'h000087F4: begin
				q			<=			16'h0113;
		end
		32'h000087F6: begin
				q			<=			16'h0301;
		end
		32'h000087F8: begin
				q			<=			16'h8067;
		end
		32'h000087FA: begin
				q			<=			16'h0000;
		end
		32'h000087FC: begin
				q			<=			16'h0737;
		end
		32'h000087FE: begin
				q			<=			16'hFFF0;
		end
		32'h00008800: begin
				q			<=			16'h87B3;
		end
		32'h00008802: begin
				q			<=			16'h02E7;
		end
		32'h00008804: begin
				q			<=			16'h8633;
		end
		32'h00008806: begin
				q			<=			16'h00B7;
		end
		32'h00008808: begin
				q			<=			16'hF06F;
		end
		32'h0000880A: begin
				q			<=			16'hFB9F;
		end
		32'h0000880C: begin
				q			<=			16'h0113;
		end
		32'h0000880E: begin
				q			<=			16'hFF01;
		end
		32'h00008810: begin
				q			<=			16'h2423;
		end
		32'h00008812: begin
				q			<=			16'h0081;
		end
		32'h00008814: begin
				q			<=			16'h2623;
		end
		32'h00008816: begin
				q			<=			16'h0011;
		end
		32'h00008818: begin
				q			<=			16'h2223;
		end
		32'h0000881A: begin
				q			<=			16'h0121;
		end
		32'h0000881C: begin
				q			<=			16'h2023;
		end
		32'h0000881E: begin
				q			<=			16'h0131;
		end
		32'h00008820: begin
				q			<=			16'h0793;
		end
		32'h00008822: begin
				q			<=			16'h0170;
		end
		32'h00008824: begin
				q			<=			16'h0413;
		end
		32'h00008826: begin
				q			<=			16'h0005;
		end
		32'h00008828: begin
				q			<=			16'hCA63;
		end
		32'h0000882A: begin
				q			<=			16'h02A7;
		end
		32'h0000882C: begin
				q			<=			16'h1413;
		end
		32'h0000882E: begin
				q			<=			16'h0035;
		end
		32'h00008830: begin
				q			<=			16'h7797;
		end
		32'h00008832: begin
				q			<=			16'h0000;
		end
		32'h00008834: begin
				q			<=			16'h8793;
		end
		32'h00008836: begin
				q			<=			16'hCD07;
		end
		32'h00008838: begin
				q			<=			16'h8433;
		end
		32'h0000883A: begin
				q			<=			16'h0087;
		end
		32'h0000883C: begin
				q			<=			16'h2503;
		end
		32'h0000883E: begin
				q			<=			16'h0104;
		end
		32'h00008840: begin
				q			<=			16'h2583;
		end
		32'h00008842: begin
				q			<=			16'h0144;
		end
		32'h00008844: begin
				q			<=			16'h2083;
		end
		32'h00008846: begin
				q			<=			16'h00C1;
		end
		32'h00008848: begin
				q			<=			16'h2403;
		end
		32'h0000884A: begin
				q			<=			16'h0081;
		end
		32'h0000884C: begin
				q			<=			16'h2903;
		end
		32'h0000884E: begin
				q			<=			16'h0041;
		end
		32'h00008850: begin
				q			<=			16'h2983;
		end
		32'h00008852: begin
				q			<=			16'h0001;
		end
		32'h00008854: begin
				q			<=			16'h0113;
		end
		32'h00008856: begin
				q			<=			16'h0101;
		end
		32'h00008858: begin
				q			<=			16'h8067;
		end
		32'h0000885A: begin
				q			<=			16'h0000;
		end
		32'h0000885C: begin
				q			<=			16'h7797;
		end
		32'h0000885E: begin
				q			<=			16'h0000;
		end
		32'h00008860: begin
				q			<=			16'h8793;
		end
		32'h00008862: begin
				q			<=			16'h6C47;
		end
		32'h00008864: begin
				q			<=			16'hA503;
		end
		32'h00008866: begin
				q			<=			16'h0007;
		end
		32'h00008868: begin
				q			<=			16'hA583;
		end
		32'h0000886A: begin
				q			<=			16'h0047;
		end
		32'h0000886C: begin
				q			<=			16'h7797;
		end
		32'h0000886E: begin
				q			<=			16'h0000;
		end
		32'h00008870: begin
				q			<=			16'h8793;
		end
		32'h00008872: begin
				q			<=			16'h6BC7;
		end
		32'h00008874: begin
				q			<=			16'hA903;
		end
		32'h00008876: begin
				q			<=			16'h0007;
		end
		32'h00008878: begin
				q			<=			16'hA983;
		end
		32'h0000887A: begin
				q			<=			16'h0047;
		end
		32'h0000887C: begin
				q			<=			16'h0613;
		end
		32'h0000887E: begin
				q			<=			16'h0009;
		end
		32'h00008880: begin
				q			<=			16'h8693;
		end
		32'h00008882: begin
				q			<=			16'h0009;
		end
		32'h00008884: begin
				q			<=			16'h0413;
		end
		32'h00008886: begin
				q			<=			16'hFFF4;
		end
		32'h00008888: begin
				q			<=			16'h30EF;
		end
		32'h0000888A: begin
				q			<=			16'h1540;
		end
		32'h0000888C: begin
				q			<=			16'h18E3;
		end
		32'h0000888E: begin
				q			<=			16'hFE04;
		end
		32'h00008890: begin
				q			<=			16'hF06F;
		end
		32'h00008892: begin
				q			<=			16'hFB5F;
		end
		32'h00008894: begin
				q			<=			16'h8793;
		end
		32'h00008896: begin
				q			<=			16'hFFF5;
		end
		32'h00008898: begin
				q			<=			16'h2703;
		end
		32'h0000889A: begin
				q			<=			16'h0106;
		end
		32'h0000889C: begin
				q			<=			16'hD793;
		end
		32'h0000889E: begin
				q			<=			16'h4057;
		end
		32'h000088A0: begin
				q			<=			16'h8793;
		end
		32'h000088A2: begin
				q			<=			16'h0017;
		end
		32'h000088A4: begin
				q			<=			16'h9793;
		end
		32'h000088A6: begin
				q			<=			16'h0027;
		end
		32'h000088A8: begin
				q			<=			16'h0693;
		end
		32'h000088AA: begin
				q			<=			16'h0146;
		end
		32'h000088AC: begin
				q			<=			16'h1713;
		end
		32'h000088AE: begin
				q			<=			16'h0027;
		end
		32'h000088B0: begin
				q			<=			16'h07B3;
		end
		32'h000088B2: begin
				q			<=			16'h00F5;
		end
		32'h000088B4: begin
				q			<=			16'h8733;
		end
		32'h000088B6: begin
				q			<=			16'h00E6;
		end
		32'h000088B8: begin
				q			<=			16'hE663;
		end
		32'h000088BA: begin
				q			<=			16'h00E6;
		end
		32'h000088BC: begin
				q			<=			16'h6E63;
		end
		32'h000088BE: begin
				q			<=			16'h00F5;
		end
		32'h000088C0: begin
				q			<=			16'h8067;
		end
		32'h000088C2: begin
				q			<=			16'h0000;
		end
		32'h000088C4: begin
				q			<=			16'h8693;
		end
		32'h000088C6: begin
				q			<=			16'h0046;
		end
		32'h000088C8: begin
				q			<=			16'hA603;
		end
		32'h000088CA: begin
				q			<=			16'hFFC6;
		end
		32'h000088CC: begin
				q			<=			16'h0513;
		end
		32'h000088CE: begin
				q			<=			16'h0045;
		end
		32'h000088D0: begin
				q			<=			16'h2E23;
		end
		32'h000088D2: begin
				q			<=			16'hFEC5;
		end
		32'h000088D4: begin
				q			<=			16'hF06F;
		end
		32'h000088D6: begin
				q			<=			16'hFE5F;
		end
		32'h000088D8: begin
				q			<=			16'h0513;
		end
		32'h000088DA: begin
				q			<=			16'h0045;
		end
		32'h000088DC: begin
				q			<=			16'h2E23;
		end
		32'h000088DE: begin
				q			<=			16'hFE05;
		end
		32'h000088E0: begin
				q			<=			16'hF06F;
		end
		32'h000088E2: begin
				q			<=			16'hFDDF;
		end
		32'h000088E4: begin
				q			<=			16'h2683;
		end
		32'h000088E6: begin
				q			<=			16'h0105;
		end
		32'h000088E8: begin
				q			<=			16'hD793;
		end
		32'h000088EA: begin
				q			<=			16'h4055;
		end
		32'h000088EC: begin
				q			<=			16'h0713;
		end
		32'h000088EE: begin
				q			<=			16'h0145;
		end
		32'h000088F0: begin
				q			<=			16'hC063;
		end
		32'h000088F2: begin
				q			<=			16'h04F6;
		end
		32'h000088F4: begin
				q			<=			16'hD463;
		end
		32'h000088F6: begin
				q			<=			16'h02D7;
		end
		32'h000088F8: begin
				q			<=			16'hF593;
		end
		32'h000088FA: begin
				q			<=			16'h01F5;
		end
		32'h000088FC: begin
				q			<=			16'h8063;
		end
		32'h000088FE: begin
				q			<=			16'h0205;
		end
		32'h00008900: begin
				q			<=			16'h9693;
		end
		32'h00008902: begin
				q			<=			16'h0027;
		end
		32'h00008904: begin
				q			<=			16'h06B3;
		end
		32'h00008906: begin
				q			<=			16'h00D7;
		end
		32'h00008908: begin
				q			<=			16'hA603;
		end
		32'h0000890A: begin
				q			<=			16'h0006;
		end
		32'h0000890C: begin
				q			<=			16'h0513;
		end
		32'h0000890E: begin
				q			<=			16'h0010;
		end
		32'h00008910: begin
				q			<=			16'h56B3;
		end
		32'h00008912: begin
				q			<=			16'h00B6;
		end
		32'h00008914: begin
				q			<=			16'h95B3;
		end
		32'h00008916: begin
				q			<=			16'h00B6;
		end
		32'h00008918: begin
				q			<=			16'h1863;
		end
		32'h0000891A: begin
				q			<=			16'h02B6;
		end
		32'h0000891C: begin
				q			<=			16'h9793;
		end
		32'h0000891E: begin
				q			<=			16'h0027;
		end
		32'h00008920: begin
				q			<=			16'h07B3;
		end
		32'h00008922: begin
				q			<=			16'h00F7;
		end
		32'h00008924: begin
				q			<=			16'h6A63;
		end
		32'h00008926: begin
				q			<=			16'h00F7;
		end
		32'h00008928: begin
				q			<=			16'h0513;
		end
		32'h0000892A: begin
				q			<=			16'h0000;
		end
		32'h0000892C: begin
				q			<=			16'h8067;
		end
		32'h0000892E: begin
				q			<=			16'h0000;
		end
		32'h00008930: begin
				q			<=			16'h8793;
		end
		32'h00008932: begin
				q			<=			16'h0006;
		end
		32'h00008934: begin
				q			<=			16'hF06F;
		end
		32'h00008936: begin
				q			<=			16'hFE9F;
		end
		32'h00008938: begin
				q			<=			16'h8793;
		end
		32'h0000893A: begin
				q			<=			16'hFFC7;
		end
		32'h0000893C: begin
				q			<=			16'hA683;
		end
		32'h0000893E: begin
				q			<=			16'h0007;
		end
		32'h00008940: begin
				q			<=			16'h82E3;
		end
		32'h00008942: begin
				q			<=			16'hFE06;
		end
		32'h00008944: begin
				q			<=			16'h0513;
		end
		32'h00008946: begin
				q			<=			16'h0010;
		end
		32'h00008948: begin
				q			<=			16'h8067;
		end
		32'h0000894A: begin
				q			<=			16'h0000;
		end
		32'h0000894C: begin
				q			<=			16'h0000;
		end
		32'h0000894E: begin
				q			<=			16'h0000;
		end
		32'h00008950: begin
				q			<=			16'h0113;
		end
		32'h00008952: begin
				q			<=			16'hFF01;
		end
		32'h00008954: begin
				q			<=			16'h2223;
		end
		32'h00008956: begin
				q			<=			16'h0091;
		end
		32'h00008958: begin
				q			<=			16'h04B7;
		end
		32'h0000895A: begin
				q			<=			16'h8000;
		end
		32'h0000895C: begin
				q			<=			16'h2423;
		end
		32'h0000895E: begin
				q			<=			16'h0081;
		end
		32'h00008960: begin
				q			<=			16'h2623;
		end
		32'h00008962: begin
				q			<=			16'h0011;
		end
		32'h00008964: begin
				q			<=			16'hC493;
		end
		32'h00008966: begin
				q			<=			16'hFFF4;
		end
		32'h00008968: begin
				q			<=			16'hF733;
		end
		32'h0000896A: begin
				q			<=			16'h00B4;
		end
		32'h0000896C: begin
				q			<=			16'h2023;
		end
		32'h0000896E: begin
				q			<=			16'h0006;
		end
		32'h00008970: begin
				q			<=			16'h0837;
		end
		32'h00008972: begin
				q			<=			16'h7FF0;
		end
		32'h00008974: begin
				q			<=			16'h0693;
		end
		32'h00008976: begin
				q			<=			16'h0005;
		end
		32'h00008978: begin
				q			<=			16'h8793;
		end
		32'h0000897A: begin
				q			<=			16'h0005;
		end
		32'h0000897C: begin
				q			<=			16'h0413;
		end
		32'h0000897E: begin
				q			<=			16'h0006;
		end
		32'h00008980: begin
				q			<=			16'h5463;
		end
		32'h00008982: begin
				q			<=			16'h0707;
		end
		32'h00008984: begin
				q			<=			16'h6833;
		end
		32'h00008986: begin
				q			<=			16'h00A7;
		end
		32'h00008988: begin
				q			<=			16'h0063;
		end
		32'h0000898A: begin
				q			<=			16'h0608;
		end
		32'h0000898C: begin
				q			<=			16'h07B7;
		end
		32'h0000898E: begin
				q			<=			16'h0010;
		end
		32'h00008990: begin
				q			<=			16'h8613;
		end
		32'h00008992: begin
				q			<=			16'h0005;
		end
		32'h00008994: begin
				q			<=			16'h5663;
		end
		32'h00008996: begin
				q			<=			16'h02F7;
		end
		32'h00008998: begin
				q			<=			16'h7797;
		end
		32'h0000899A: begin
				q			<=			16'h0000;
		end
		32'h0000899C: begin
				q			<=			16'h8793;
		end
		32'h0000899E: begin
				q			<=			16'h5987;
		end
		32'h000089A0: begin
				q			<=			16'hA603;
		end
		32'h000089A2: begin
				q			<=			16'h0007;
		end
		32'h000089A4: begin
				q			<=			16'hA683;
		end
		32'h000089A6: begin
				q			<=			16'h0047;
		end
		32'h000089A8: begin
				q			<=			16'h30EF;
		end
		32'h000089AA: begin
				q			<=			16'h0340;
		end
		32'h000089AC: begin
				q			<=			16'h0793;
		end
		32'h000089AE: begin
				q			<=			16'hFCA0;
		end
		32'h000089B0: begin
				q			<=			16'h0693;
		end
		32'h000089B2: begin
				q			<=			16'h0005;
		end
		32'h000089B4: begin
				q			<=			16'h8613;
		end
		32'h000089B6: begin
				q			<=			16'h0005;
		end
		32'h000089B8: begin
				q			<=			16'hF733;
		end
		32'h000089BA: begin
				q			<=			16'h00B4;
		end
		32'h000089BC: begin
				q			<=			16'h2023;
		end
		32'h000089BE: begin
				q			<=			16'h00F4;
		end
		32'h000089C0: begin
				q			<=			16'h2783;
		end
		32'h000089C2: begin
				q			<=			16'h0004;
		end
		32'h000089C4: begin
				q			<=			16'h5713;
		end
		32'h000089C6: begin
				q			<=			16'h4147;
		end
		32'h000089C8: begin
				q			<=			16'h0713;
		end
		32'h000089CA: begin
				q			<=			16'hC027;
		end
		32'h000089CC: begin
				q			<=			16'h8733;
		end
		32'h000089CE: begin
				q			<=			16'h00E7;
		end
		32'h000089D0: begin
				q			<=			16'h07B7;
		end
		32'h000089D2: begin
				q			<=			16'h8010;
		end
		32'h000089D4: begin
				q			<=			16'h8793;
		end
		32'h000089D6: begin
				q			<=			16'hFFF7;
		end
		32'h000089D8: begin
				q			<=			16'h7633;
		end
		32'h000089DA: begin
				q			<=			16'h00F6;
		end
		32'h000089DC: begin
				q			<=			16'h07B7;
		end
		32'h000089DE: begin
				q			<=			16'h3FE0;
		end
		32'h000089E0: begin
				q			<=			16'h2023;
		end
		32'h000089E2: begin
				q			<=			16'h00E4;
		end
		32'h000089E4: begin
				q			<=			16'h67B3;
		end
		32'h000089E6: begin
				q			<=			16'h00F6;
		end
		32'h000089E8: begin
				q			<=			16'h2083;
		end
		32'h000089EA: begin
				q			<=			16'h00C1;
		end
		32'h000089EC: begin
				q			<=			16'h2403;
		end
		32'h000089EE: begin
				q			<=			16'h0081;
		end
		32'h000089F0: begin
				q			<=			16'h2483;
		end
		32'h000089F2: begin
				q			<=			16'h0041;
		end
		32'h000089F4: begin
				q			<=			16'h8513;
		end
		32'h000089F6: begin
				q			<=			16'h0006;
		end
		32'h000089F8: begin
				q			<=			16'h8593;
		end
		32'h000089FA: begin
				q			<=			16'h0007;
		end
		32'h000089FC: begin
				q			<=			16'h0113;
		end
		32'h000089FE: begin
				q			<=			16'h0101;
		end
		32'h00008A00: begin
				q			<=			16'h8067;
		end
		32'h00008A02: begin
				q			<=			16'h0000;
		end
		32'h00008A04: begin
				q			<=			16'h0000;
		end
		32'h00008A06: begin
				q			<=			16'h0000;
		end
		32'h00008A08: begin
				q			<=			16'h0113;
		end
		32'h00008A0A: begin
				q			<=			16'hFF01;
		end
		32'h00008A0C: begin
				q			<=			16'h2423;
		end
		32'h00008A0E: begin
				q			<=			16'h0081;
		end
		32'h00008A10: begin
				q			<=			16'h0413;
		end
		32'h00008A12: begin
				q			<=			16'h0005;
		end
		32'h00008A14: begin
				q			<=			16'h8513;
		end
		32'h00008A16: begin
				q			<=			16'h0005;
		end
		32'h00008A18: begin
				q			<=			16'h8797;
		end
		32'h00008A1A: begin
				q			<=			16'h0000;
		end
		32'h00008A1C: begin
				q			<=			16'hAA23;
		end
		32'h00008A1E: begin
				q			<=			16'h5407;
		end
		32'h00008A20: begin
				q			<=			16'h2623;
		end
		32'h00008A22: begin
				q			<=			16'h0011;
		end
		32'h00008A24: begin
				q			<=			16'h10EF;
		end
		32'h00008A26: begin
				q			<=			16'h7AD0;
		end
		32'h00008A28: begin
				q			<=			16'h0793;
		end
		32'h00008A2A: begin
				q			<=			16'hFFF0;
		end
		32'h00008A2C: begin
				q			<=			16'h1C63;
		end
		32'h00008A2E: begin
				q			<=			16'h00F5;
		end
		32'h00008A30: begin
				q			<=			16'h8797;
		end
		32'h00008A32: begin
				q			<=			16'h0000;
		end
		32'h00008A34: begin
				q			<=			16'h8793;
		end
		32'h00008A36: begin
				q			<=			16'h53C7;
		end
		32'h00008A38: begin
				q			<=			16'hA783;
		end
		32'h00008A3A: begin
				q			<=			16'h0007;
		end
		32'h00008A3C: begin
				q			<=			16'h8463;
		end
		32'h00008A3E: begin
				q			<=			16'h0007;
		end
		32'h00008A40: begin
				q			<=			16'h2023;
		end
		32'h00008A42: begin
				q			<=			16'h00F4;
		end
		32'h00008A44: begin
				q			<=			16'h2083;
		end
		32'h00008A46: begin
				q			<=			16'h00C1;
		end
		32'h00008A48: begin
				q			<=			16'h2403;
		end
		32'h00008A4A: begin
				q			<=			16'h0081;
		end
		32'h00008A4C: begin
				q			<=			16'h0113;
		end
		32'h00008A4E: begin
				q			<=			16'h0101;
		end
		32'h00008A50: begin
				q			<=			16'h8067;
		end
		32'h00008A52: begin
				q			<=			16'h0000;
		end
		32'h00008A54: begin
				q			<=			16'h0000;
		end
		32'h00008A56: begin
				q			<=			16'h0000;
		end
		32'h00008A58: begin
				q			<=			16'h0113;
		end
		32'h00008A5A: begin
				q			<=			16'hF601;
		end
		32'h00008A5C: begin
				q			<=			16'h2A23;
		end
		32'h00008A5E: begin
				q			<=			16'h08F1;
		end
		32'h00008A60: begin
				q			<=			16'h07B7;
		end
		32'h00008A62: begin
				q			<=			16'h8000;
		end
		32'h00008A64: begin
				q			<=			16'hC793;
		end
		32'h00008A66: begin
				q			<=			16'hFFF7;
		end
		32'h00008A68: begin
				q			<=			16'h2E23;
		end
		32'h00008A6A: begin
				q			<=			16'h00F1;
		end
		32'h00008A6C: begin
				q			<=			16'h2823;
		end
		32'h00008A6E: begin
				q			<=			16'h00F1;
		end
		32'h00008A70: begin
				q			<=			16'h07B7;
		end
		32'h00008A72: begin
				q			<=			16'hFFFF;
		end
		32'h00008A74: begin
				q			<=			16'h2623;
		end
		32'h00008A76: begin
				q			<=			16'h08D1;
		end
		32'h00008A78: begin
				q			<=			16'h2423;
		end
		32'h00008A7A: begin
				q			<=			16'h00B1;
		end
		32'h00008A7C: begin
				q			<=			16'h2C23;
		end
		32'h00008A7E: begin
				q			<=			16'h00B1;
		end
		32'h00008A80: begin
				q			<=			16'h8793;
		end
		32'h00008A82: begin
				q			<=			16'h2087;
		end
		32'h00008A84: begin
				q			<=			16'h0693;
		end
		32'h00008A86: begin
				q			<=			16'h08C1;
		end
		32'h00008A88: begin
				q			<=			16'h0593;
		end
		32'h00008A8A: begin
				q			<=			16'h0081;
		end
		32'h00008A8C: begin
				q			<=			16'h2E23;
		end
		32'h00008A8E: begin
				q			<=			16'h0611;
		end
		32'h00008A90: begin
				q			<=			16'h2A23;
		end
		32'h00008A92: begin
				q			<=			16'h00F1;
		end
		32'h00008A94: begin
				q			<=			16'h2823;
		end
		32'h00008A96: begin
				q			<=			16'h08E1;
		end
		32'h00008A98: begin
				q			<=			16'h2C23;
		end
		32'h00008A9A: begin
				q			<=			16'h0901;
		end
		32'h00008A9C: begin
				q			<=			16'h2E23;
		end
		32'h00008A9E: begin
				q			<=			16'h0911;
		end
		32'h00008AA0: begin
				q			<=			16'h2223;
		end
		32'h00008AA2: begin
				q			<=			16'h00D1;
		end
		32'h00008AA4: begin
				q			<=			16'hA0EF;
		end
		32'h00008AA6: begin
				q			<=			16'hC34F;
		end
		32'h00008AA8: begin
				q			<=			16'h2783;
		end
		32'h00008AAA: begin
				q			<=			16'h0081;
		end
		32'h00008AAC: begin
				q			<=			16'h8023;
		end
		32'h00008AAE: begin
				q			<=			16'h0007;
		end
		32'h00008AB0: begin
				q			<=			16'h2083;
		end
		32'h00008AB2: begin
				q			<=			16'h07C1;
		end
		32'h00008AB4: begin
				q			<=			16'h0113;
		end
		32'h00008AB6: begin
				q			<=			16'h0A01;
		end
		32'h00008AB8: begin
				q			<=			16'h8067;
		end
		32'h00008ABA: begin
				q			<=			16'h0000;
		end
		32'h00008ABC: begin
				q			<=			16'h0113;
		end
		32'h00008ABE: begin
				q			<=			16'hF601;
		end
		32'h00008AC0: begin
				q			<=			16'h2A23;
		end
		32'h00008AC2: begin
				q			<=			16'h08F1;
		end
		32'h00008AC4: begin
				q			<=			16'h07B7;
		end
		32'h00008AC6: begin
				q			<=			16'h8000;
		end
		32'h00008AC8: begin
				q			<=			16'hC793;
		end
		32'h00008ACA: begin
				q			<=			16'hFFF7;
		end
		32'h00008ACC: begin
				q			<=			16'h2E23;
		end
		32'h00008ACE: begin
				q			<=			16'h00F1;
		end
		32'h00008AD0: begin
				q			<=			16'h2823;
		end
		32'h00008AD2: begin
				q			<=			16'h00F1;
		end
		32'h00008AD4: begin
				q			<=			16'h07B7;
		end
		32'h00008AD6: begin
				q			<=			16'hFFFF;
		end
		32'h00008AD8: begin
				q			<=			16'h8793;
		end
		32'h00008ADA: begin
				q			<=			16'h2087;
		end
		32'h00008ADC: begin
				q			<=			16'h2423;
		end
		32'h00008ADE: begin
				q			<=			16'h08C1;
		end
		32'h00008AE0: begin
				q			<=			16'h2623;
		end
		32'h00008AE2: begin
				q			<=			16'h08D1;
		end
		32'h00008AE4: begin
				q			<=			16'h2823;
		end
		32'h00008AE6: begin
				q			<=			16'h08E1;
		end
		32'h00008AE8: begin
				q			<=			16'h2C23;
		end
		32'h00008AEA: begin
				q			<=			16'h0901;
		end
		32'h00008AEC: begin
				q			<=			16'h2E23;
		end
		32'h00008AEE: begin
				q			<=			16'h0911;
		end
		32'h00008AF0: begin
				q			<=			16'h2A23;
		end
		32'h00008AF2: begin
				q			<=			16'h00F1;
		end
		32'h00008AF4: begin
				q			<=			16'h8797;
		end
		32'h00008AF6: begin
				q			<=			16'h0000;
		end
		32'h00008AF8: begin
				q			<=			16'h8793;
		end
		32'h00008AFA: begin
				q			<=			16'hDE47;
		end
		32'h00008AFC: begin
				q			<=			16'h2423;
		end
		32'h00008AFE: begin
				q			<=			16'h00A1;
		end
		32'h00008B00: begin
				q			<=			16'h2C23;
		end
		32'h00008B02: begin
				q			<=			16'h00A1;
		end
		32'h00008B04: begin
				q			<=			16'hA503;
		end
		32'h00008B06: begin
				q			<=			16'h0007;
		end
		32'h00008B08: begin
				q			<=			16'h0693;
		end
		32'h00008B0A: begin
				q			<=			16'h0881;
		end
		32'h00008B0C: begin
				q			<=			16'h8613;
		end
		32'h00008B0E: begin
				q			<=			16'h0005;
		end
		32'h00008B10: begin
				q			<=			16'h0593;
		end
		32'h00008B12: begin
				q			<=			16'h0081;
		end
		32'h00008B14: begin
				q			<=			16'h2E23;
		end
		32'h00008B16: begin
				q			<=			16'h0611;
		end
		32'h00008B18: begin
				q			<=			16'h2223;
		end
		32'h00008B1A: begin
				q			<=			16'h00D1;
		end
		32'h00008B1C: begin
				q			<=			16'hA097;
		end
		32'h00008B1E: begin
				q			<=			16'hFFFF;
		end
		32'h00008B20: begin
				q			<=			16'h80E7;
		end
		32'h00008B22: begin
				q			<=			16'h3BC0;
		end
		32'h00008B24: begin
				q			<=			16'h2783;
		end
		32'h00008B26: begin
				q			<=			16'h0081;
		end
		32'h00008B28: begin
				q			<=			16'h8023;
		end
		32'h00008B2A: begin
				q			<=			16'h0007;
		end
		32'h00008B2C: begin
				q			<=			16'h2083;
		end
		32'h00008B2E: begin
				q			<=			16'h07C1;
		end
		32'h00008B30: begin
				q			<=			16'h0113;
		end
		32'h00008B32: begin
				q			<=			16'h0A01;
		end
		32'h00008B34: begin
				q			<=			16'h8067;
		end
		32'h00008B36: begin
				q			<=			16'h0000;
		end
		32'h00008B38: begin
				q			<=			16'h0000;
		end
		32'h00008B3A: begin
				q			<=			16'h0000;
		end
		32'h00008B3C: begin
				q			<=			16'h0793;
		end
		32'h00008B3E: begin
				q			<=			16'h0005;
		end
		32'h00008B40: begin
				q			<=			16'hC703;
		end
		32'h00008B42: begin
				q			<=			16'h0005;
		end
		32'h00008B44: begin
				q			<=			16'h8793;
		end
		32'h00008B46: begin
				q			<=			16'h0017;
		end
		32'h00008B48: begin
				q			<=			16'h8593;
		end
		32'h00008B4A: begin
				q			<=			16'h0015;
		end
		32'h00008B4C: begin
				q			<=			16'h8FA3;
		end
		32'h00008B4E: begin
				q			<=			16'hFEE7;
		end
		32'h00008B50: begin
				q			<=			16'h18E3;
		end
		32'h00008B52: begin
				q			<=			16'hFE07;
		end
		32'h00008B54: begin
				q			<=			16'h8067;
		end
		32'h00008B56: begin
				q			<=			16'h0000;
		end
		32'h00008B58: begin
				q			<=			16'h0000;
		end
		32'h00008B5A: begin
				q			<=			16'h0000;
		end
		32'h00008B5C: begin
				q			<=			16'h2783;
		end
		32'h00008B5E: begin
				q			<=			16'h0086;
		end
		32'h00008B60: begin
				q			<=			16'h0113;
		end
		32'h00008B62: begin
				q			<=			16'hFD01;
		end
		32'h00008B64: begin
				q			<=			16'h2E23;
		end
		32'h00008B66: begin
				q			<=			16'h0131;
		end
		32'h00008B68: begin
				q			<=			16'h2623;
		end
		32'h00008B6A: begin
				q			<=			16'h0211;
		end
		32'h00008B6C: begin
				q			<=			16'h2423;
		end
		32'h00008B6E: begin
				q			<=			16'h0281;
		end
		32'h00008B70: begin
				q			<=			16'h2223;
		end
		32'h00008B72: begin
				q			<=			16'h0291;
		end
		32'h00008B74: begin
				q			<=			16'h2023;
		end
		32'h00008B76: begin
				q			<=			16'h0321;
		end
		32'h00008B78: begin
				q			<=			16'h2C23;
		end
		32'h00008B7A: begin
				q			<=			16'h0141;
		end
		32'h00008B7C: begin
				q			<=			16'h2A23;
		end
		32'h00008B7E: begin
				q			<=			16'h0151;
		end
		32'h00008B80: begin
				q			<=			16'h2823;
		end
		32'h00008B82: begin
				q			<=			16'h0161;
		end
		32'h00008B84: begin
				q			<=			16'h2623;
		end
		32'h00008B86: begin
				q			<=			16'h0171;
		end
		32'h00008B88: begin
				q			<=			16'h2423;
		end
		32'h00008B8A: begin
				q			<=			16'h0181;
		end
		32'h00008B8C: begin
				q			<=			16'h2223;
		end
		32'h00008B8E: begin
				q			<=			16'h0191;
		end
		32'h00008B90: begin
				q			<=			16'h2023;
		end
		32'h00008B92: begin
				q			<=			16'h01A1;
		end
		32'h00008B94: begin
				q			<=			16'h0993;
		end
		32'h00008B96: begin
				q			<=			16'h0006;
		end
		32'h00008B98: begin
				q			<=			16'h8463;
		end
		32'h00008B9A: begin
				q			<=			16'h1207;
		end
		32'h00008B9C: begin
				q			<=			16'h2A83;
		end
		32'h00008B9E: begin
				q			<=			16'h0006;
		end
		32'h00008BA0: begin
				q			<=			16'h0A13;
		end
		32'h00008BA2: begin
				q			<=			16'h0005;
		end
		32'h00008BA4: begin
				q			<=			16'h8413;
		end
		32'h00008BA6: begin
				q			<=			16'h0005;
		end
		32'h00008BA8: begin
				q			<=			16'h0B13;
		end
		32'h00008BAA: begin
				q			<=			16'h0000;
		end
		32'h00008BAC: begin
				q			<=			16'h0913;
		end
		32'h00008BAE: begin
				q			<=			16'h0000;
		end
		32'h00008BB0: begin
				q			<=			16'h0B93;
		end
		32'h00008BB2: begin
				q			<=			16'h0030;
		end
		32'h00008BB4: begin
				q			<=			16'h0C13;
		end
		32'h00008BB6: begin
				q			<=			16'h0020;
		end
		32'h00008BB8: begin
				q			<=			16'h0063;
		end
		32'h00008BBA: begin
				q			<=			16'h0809;
		end
		32'h00008BBC: begin
				q			<=			16'h2D03;
		end
		32'h00008BBE: begin
				q			<=			16'h0084;
		end
		32'h00008BC0: begin
				q			<=			16'h6063;
		end
		32'h00008BC2: begin
				q			<=			16'h0DA9;
		end
		32'h00008BC4: begin
				q			<=			16'h5783;
		end
		32'h00008BC6: begin
				q			<=			16'h00C4;
		end
		32'h00008BC8: begin
				q			<=			16'hF713;
		end
		32'h00008BCA: begin
				q			<=			16'h4807;
		end
		32'h00008BCC: begin
				q			<=			16'h0A63;
		end
		32'h00008BCE: begin
				q			<=			16'h0A07;
		end
		32'h00008BD0: begin
				q			<=			16'h2483;
		end
		32'h00008BD2: begin
				q			<=			16'h0004;
		end
		32'h00008BD4: begin
				q			<=			16'h2583;
		end
		32'h00008BD6: begin
				q			<=			16'h0104;
		end
		32'h00008BD8: begin
				q			<=			16'h8CB3;
		end
		32'h00008BDA: begin
				q			<=			16'h40B4;
		end
		32'h00008BDC: begin
				q			<=			16'h2483;
		end
		32'h00008BDE: begin
				q			<=			16'h0144;
		end
		32'h00008BE0: begin
				q			<=			16'h8713;
		end
		32'h00008BE2: begin
				q			<=			16'h001C;
		end
		32'h00008BE4: begin
				q			<=			16'h0733;
		end
		32'h00008BE6: begin
				q			<=			16'h0127;
		end
		32'h00008BE8: begin
				q			<=			16'h84B3;
		end
		32'h00008BEA: begin
				q			<=			16'h029B;
		end
		32'h00008BEC: begin
				q			<=			16'hC4B3;
		end
		32'h00008BEE: begin
				q			<=			16'h0384;
		end
		32'h00008BF0: begin
				q			<=			16'hF463;
		end
		32'h00008BF2: begin
				q			<=			16'h00E4;
		end
		32'h00008BF4: begin
				q			<=			16'h0493;
		end
		32'h00008BF6: begin
				q			<=			16'h0007;
		end
		32'h00008BF8: begin
				q			<=			16'hF793;
		end
		32'h00008BFA: begin
				q			<=			16'h4007;
		end
		32'h00008BFC: begin
				q			<=			16'h8263;
		end
		32'h00008BFE: begin
				q			<=			16'h1007;
		end
		32'h00008C00: begin
				q			<=			16'h8593;
		end
		32'h00008C02: begin
				q			<=			16'h0004;
		end
		32'h00008C04: begin
				q			<=			16'h0513;
		end
		32'h00008C06: begin
				q			<=			16'h000A;
		end
		32'h00008C08: begin
				q			<=			16'hE0EF;
		end
		32'h00008C0A: begin
				q			<=			16'hF98F;
		end
		32'h00008C0C: begin
				q			<=			16'h0D13;
		end
		32'h00008C0E: begin
				q			<=			16'h0005;
		end
		32'h00008C10: begin
				q			<=			16'h1C63;
		end
		32'h00008C12: begin
				q			<=			16'h0205;
		end
		32'h00008C14: begin
				q			<=			16'h0793;
		end
		32'h00008C16: begin
				q			<=			16'h00C0;
		end
		32'h00008C18: begin
				q			<=			16'h2023;
		end
		32'h00008C1A: begin
				q			<=			16'h00FA;
		end
		32'h00008C1C: begin
				q			<=			16'h5783;
		end
		32'h00008C1E: begin
				q			<=			16'h00C4;
		end
		32'h00008C20: begin
				q			<=			16'h0513;
		end
		32'h00008C22: begin
				q			<=			16'hFFF0;
		end
		32'h00008C24: begin
				q			<=			16'hE793;
		end
		32'h00008C26: begin
				q			<=			16'h0407;
		end
		32'h00008C28: begin
				q			<=			16'h1623;
		end
		32'h00008C2A: begin
				q			<=			16'h00F4;
		end
		32'h00008C2C: begin
				q			<=			16'hA423;
		end
		32'h00008C2E: begin
				q			<=			16'h0009;
		end
		32'h00008C30: begin
				q			<=			16'hA223;
		end
		32'h00008C32: begin
				q			<=			16'h0009;
		end
		32'h00008C34: begin
				q			<=			16'h006F;
		end
		32'h00008C36: begin
				q			<=			16'h0940;
		end
		32'h00008C38: begin
				q			<=			16'hAB03;
		end
		32'h00008C3A: begin
				q			<=			16'h000A;
		end
		32'h00008C3C: begin
				q			<=			16'hA903;
		end
		32'h00008C3E: begin
				q			<=			16'h004A;
		end
		32'h00008C40: begin
				q			<=			16'h8A93;
		end
		32'h00008C42: begin
				q			<=			16'h008A;
		end
		32'h00008C44: begin
				q			<=			16'hF06F;
		end
		32'h00008C46: begin
				q			<=			16'hF75F;
		end
		32'h00008C48: begin
				q			<=			16'h2583;
		end
		32'h00008C4A: begin
				q			<=			16'h0104;
		end
		32'h00008C4C: begin
				q			<=			16'h8613;
		end
		32'h00008C4E: begin
				q			<=			16'h000C;
		end
		32'h00008C50: begin
				q			<=			16'h90EF;
		end
		32'h00008C52: begin
				q			<=			16'hEA9F;
		end
		32'h00008C54: begin
				q			<=			16'h5783;
		end
		32'h00008C56: begin
				q			<=			16'h00C4;
		end
		32'h00008C58: begin
				q			<=			16'hF793;
		end
		32'h00008C5A: begin
				q			<=			16'hB7F7;
		end
		32'h00008C5C: begin
				q			<=			16'hE793;
		end
		32'h00008C5E: begin
				q			<=			16'h0807;
		end
		32'h00008C60: begin
				q			<=			16'h1623;
		end
		32'h00008C62: begin
				q			<=			16'h00F4;
		end
		32'h00008C64: begin
				q			<=			16'h2823;
		end
		32'h00008C66: begin
				q			<=			16'h01A4;
		end
		32'h00008C68: begin
				q			<=			16'h2A23;
		end
		32'h00008C6A: begin
				q			<=			16'h0094;
		end
		32'h00008C6C: begin
				q			<=			16'h0D33;
		end
		32'h00008C6E: begin
				q			<=			16'h019D;
		end
		32'h00008C70: begin
				q			<=			16'h84B3;
		end
		32'h00008C72: begin
				q			<=			16'h4194;
		end
		32'h00008C74: begin
				q			<=			16'h2023;
		end
		32'h00008C76: begin
				q			<=			16'h01A4;
		end
		32'h00008C78: begin
				q			<=			16'h2423;
		end
		32'h00008C7A: begin
				q			<=			16'h0094;
		end
		32'h00008C7C: begin
				q			<=			16'h0D13;
		end
		32'h00008C7E: begin
				q			<=			16'h0009;
		end
		32'h00008C80: begin
				q			<=			16'h7463;
		end
		32'h00008C82: begin
				q			<=			16'h01A9;
		end
		32'h00008C84: begin
				q			<=			16'h0D13;
		end
		32'h00008C86: begin
				q			<=			16'h0009;
		end
		32'h00008C88: begin
				q			<=			16'h2503;
		end
		32'h00008C8A: begin
				q			<=			16'h0004;
		end
		32'h00008C8C: begin
				q			<=			16'h0613;
		end
		32'h00008C8E: begin
				q			<=			16'h000D;
		end
		32'h00008C90: begin
				q			<=			16'h0593;
		end
		32'h00008C92: begin
				q			<=			16'h000B;
		end
		32'h00008C94: begin
				q			<=			16'h00EF;
		end
		32'h00008C96: begin
				q			<=			16'h7490;
		end
		32'h00008C98: begin
				q			<=			16'h2783;
		end
		32'h00008C9A: begin
				q			<=			16'h0084;
		end
		32'h00008C9C: begin
				q			<=			16'h87B3;
		end
		32'h00008C9E: begin
				q			<=			16'h41A7;
		end
		32'h00008CA0: begin
				q			<=			16'h2423;
		end
		32'h00008CA2: begin
				q			<=			16'h00F4;
		end
		32'h00008CA4: begin
				q			<=			16'h2783;
		end
		32'h00008CA6: begin
				q			<=			16'h0004;
		end
		32'h00008CA8: begin
				q			<=			16'h8D33;
		end
		32'h00008CAA: begin
				q			<=			16'h01A7;
		end
		32'h00008CAC: begin
				q			<=			16'hA783;
		end
		32'h00008CAE: begin
				q			<=			16'h0089;
		end
		32'h00008CB0: begin
				q			<=			16'h2023;
		end
		32'h00008CB2: begin
				q			<=			16'h01A4;
		end
		32'h00008CB4: begin
				q			<=			16'h8933;
		end
		32'h00008CB6: begin
				q			<=			16'h4127;
		end
		32'h00008CB8: begin
				q			<=			16'hA423;
		end
		32'h00008CBA: begin
				q			<=			16'h0129;
		end
		32'h00008CBC: begin
				q			<=			16'h1EE3;
		end
		32'h00008CBE: begin
				q			<=			16'hF609;
		end
		32'h00008CC0: begin
				q			<=			16'hA223;
		end
		32'h00008CC2: begin
				q			<=			16'h0009;
		end
		32'h00008CC4: begin
				q			<=			16'h0513;
		end
		32'h00008CC6: begin
				q			<=			16'h0000;
		end
		32'h00008CC8: begin
				q			<=			16'h2083;
		end
		32'h00008CCA: begin
				q			<=			16'h02C1;
		end
		32'h00008CCC: begin
				q			<=			16'h2403;
		end
		32'h00008CCE: begin
				q			<=			16'h0281;
		end
		32'h00008CD0: begin
				q			<=			16'h2483;
		end
		32'h00008CD2: begin
				q			<=			16'h0241;
		end
		32'h00008CD4: begin
				q			<=			16'h2903;
		end
		32'h00008CD6: begin
				q			<=			16'h0201;
		end
		32'h00008CD8: begin
				q			<=			16'h2983;
		end
		32'h00008CDA: begin
				q			<=			16'h01C1;
		end
		32'h00008CDC: begin
				q			<=			16'h2A03;
		end
		32'h00008CDE: begin
				q			<=			16'h0181;
		end
		32'h00008CE0: begin
				q			<=			16'h2A83;
		end
		32'h00008CE2: begin
				q			<=			16'h0141;
		end
		32'h00008CE4: begin
				q			<=			16'h2B03;
		end
		32'h00008CE6: begin
				q			<=			16'h0101;
		end
		32'h00008CE8: begin
				q			<=			16'h2B83;
		end
		32'h00008CEA: begin
				q			<=			16'h00C1;
		end
		32'h00008CEC: begin
				q			<=			16'h2C03;
		end
		32'h00008CEE: begin
				q			<=			16'h0081;
		end
		32'h00008CF0: begin
				q			<=			16'h2C83;
		end
		32'h00008CF2: begin
				q			<=			16'h0041;
		end
		32'h00008CF4: begin
				q			<=			16'h2D03;
		end
		32'h00008CF6: begin
				q			<=			16'h0001;
		end
		32'h00008CF8: begin
				q			<=			16'h0113;
		end
		32'h00008CFA: begin
				q			<=			16'h0301;
		end
		32'h00008CFC: begin
				q			<=			16'h8067;
		end
		32'h00008CFE: begin
				q			<=			16'h0000;
		end
		32'h00008D00: begin
				q			<=			16'h8613;
		end
		32'h00008D02: begin
				q			<=			16'h0004;
		end
		32'h00008D04: begin
				q			<=			16'h0513;
		end
		32'h00008D06: begin
				q			<=			16'h000A;
		end
		32'h00008D08: begin
				q			<=			16'h00EF;
		end
		32'h00008D0A: begin
				q			<=			16'h72D0;
		end
		32'h00008D0C: begin
				q			<=			16'h0D13;
		end
		32'h00008D0E: begin
				q			<=			16'h0005;
		end
		32'h00008D10: begin
				q			<=			16'h1AE3;
		end
		32'h00008D12: begin
				q			<=			16'hF405;
		end
		32'h00008D14: begin
				q			<=			16'h2583;
		end
		32'h00008D16: begin
				q			<=			16'h0104;
		end
		32'h00008D18: begin
				q			<=			16'h0513;
		end
		32'h00008D1A: begin
				q			<=			16'h000A;
		end
		32'h00008D1C: begin
				q			<=			16'hC097;
		end
		32'h00008D1E: begin
				q			<=			16'hFFFF;
		end
		32'h00008D20: begin
				q			<=			16'h80E7;
		end
		32'h00008D22: begin
				q			<=			16'h2540;
		end
		32'h00008D24: begin
				q			<=			16'hF06F;
		end
		32'h00008D26: begin
				q			<=			16'hEF1F;
		end
		32'h00008D28: begin
				q			<=			16'hD783;
		end
		32'h00008D2A: begin
				q			<=			16'h00C5;
		end
		32'h00008D2C: begin
				q			<=			16'h0113;
		end
		32'h00008D2E: begin
				q			<=			16'hED01;
		end
		32'h00008D30: begin
				q			<=			16'h2223;
		end
		32'h00008D32: begin
				q			<=			16'h1291;
		end
		32'h00008D34: begin
				q			<=			16'h2023;
		end
		32'h00008D36: begin
				q			<=			16'h1321;
		end
		32'h00008D38: begin
				q			<=			16'h2E23;
		end
		32'h00008D3A: begin
				q			<=			16'h1131;
		end
		32'h00008D3C: begin
				q			<=			16'h2A23;
		end
		32'h00008D3E: begin
				q			<=			16'h1151;
		end
		32'h00008D40: begin
				q			<=			16'h2623;
		end
		32'h00008D42: begin
				q			<=			16'h1211;
		end
		32'h00008D44: begin
				q			<=			16'h2423;
		end
		32'h00008D46: begin
				q			<=			16'h1281;
		end
		32'h00008D48: begin
				q			<=			16'h2C23;
		end
		32'h00008D4A: begin
				q			<=			16'h1141;
		end
		32'h00008D4C: begin
				q			<=			16'h2823;
		end
		32'h00008D4E: begin
				q			<=			16'h1161;
		end
		32'h00008D50: begin
				q			<=			16'h2623;
		end
		32'h00008D52: begin
				q			<=			16'h1171;
		end
		32'h00008D54: begin
				q			<=			16'h2423;
		end
		32'h00008D56: begin
				q			<=			16'h1181;
		end
		32'h00008D58: begin
				q			<=			16'h2223;
		end
		32'h00008D5A: begin
				q			<=			16'h1191;
		end
		32'h00008D5C: begin
				q			<=			16'h2023;
		end
		32'h00008D5E: begin
				q			<=			16'h11A1;
		end
		32'h00008D60: begin
				q			<=			16'h2E23;
		end
		32'h00008D62: begin
				q			<=			16'h0FB1;
		end
		32'h00008D64: begin
				q			<=			16'hF793;
		end
		32'h00008D66: begin
				q			<=			16'h0807;
		end
		32'h00008D68: begin
				q			<=			16'h0A93;
		end
		32'h00008D6A: begin
				q			<=			16'h0005;
		end
		32'h00008D6C: begin
				q			<=			16'h8913;
		end
		32'h00008D6E: begin
				q			<=			16'h0005;
		end
		32'h00008D70: begin
				q			<=			16'h0993;
		end
		32'h00008D72: begin
				q			<=			16'h0006;
		end
		32'h00008D74: begin
				q			<=			16'h8493;
		end
		32'h00008D76: begin
				q			<=			16'h0006;
		end
		32'h00008D78: begin
				q			<=			16'h8E63;
		end
		32'h00008D7A: begin
				q			<=			16'h0207;
		end
		32'h00008D7C: begin
				q			<=			16'hA783;
		end
		32'h00008D7E: begin
				q			<=			16'h0105;
		end
		32'h00008D80: begin
				q			<=			16'h9A63;
		end
		32'h00008D82: begin
				q			<=			16'h0207;
		end
		32'h00008D84: begin
				q			<=			16'h0593;
		end
		32'h00008D86: begin
				q			<=			16'h0400;
		end
		32'h00008D88: begin
				q			<=			16'hE097;
		end
		32'h00008D8A: begin
				q			<=			16'hFFFF;
		end
		32'h00008D8C: begin
				q			<=			16'h80E7;
		end
		32'h00008D8E: begin
				q			<=			16'h6180;
		end
		32'h00008D90: begin
				q			<=			16'h2023;
		end
		32'h00008D92: begin
				q			<=			16'h00A9;
		end
		32'h00008D94: begin
				q			<=			16'h2823;
		end
		32'h00008D96: begin
				q			<=			16'h00A9;
		end
		32'h00008D98: begin
				q			<=			16'h1A63;
		end
		32'h00008D9A: begin
				q			<=			16'h0005;
		end
		32'h00008D9C: begin
				q			<=			16'h0793;
		end
		32'h00008D9E: begin
				q			<=			16'h00C0;
		end
		32'h00008DA0: begin
				q			<=			16'hA023;
		end
		32'h00008DA2: begin
				q			<=			16'h00FA;
		end
		32'h00008DA4: begin
				q			<=			16'h0B93;
		end
		32'h00008DA6: begin
				q			<=			16'hFFF0;
		end
		32'h00008DA8: begin
				q			<=			16'h006F;
		end
		32'h00008DAA: begin
				q			<=			16'h3750;
		end
		32'h00008DAC: begin
				q			<=			16'h0793;
		end
		32'h00008DAE: begin
				q			<=			16'h0400;
		end
		32'h00008DB0: begin
				q			<=			16'h2A23;
		end
		32'h00008DB2: begin
				q			<=			16'h00F9;
		end
		32'h00008DB4: begin
				q			<=			16'h0B13;
		end
		32'h00008DB6: begin
				q			<=			16'h04C1;
		end
		32'h00008DB8: begin
				q			<=			16'h2023;
		end
		32'h00008DBA: begin
				q			<=			16'h0561;
		end
		32'h00008DBC: begin
				q			<=			16'h2423;
		end
		32'h00008DBE: begin
				q			<=			16'h0401;
		end
		32'h00008DC0: begin
				q			<=			16'h2223;
		end
		32'h00008DC2: begin
				q			<=			16'h0401;
		end
		32'h00008DC4: begin
				q			<=			16'h0713;
		end
		32'h00008DC6: begin
				q			<=			16'h000B;
		end
		32'h00008DC8: begin
				q			<=			16'h2A23;
		end
		32'h00008DCA: begin
				q			<=			16'h0001;
		end
		32'h00008DCC: begin
				q			<=			16'h2623;
		end
		32'h00008DCE: begin
				q			<=			16'h0001;
		end
		32'h00008DD0: begin
				q			<=			16'h2823;
		end
		32'h00008DD2: begin
				q			<=			16'h0001;
		end
		32'h00008DD4: begin
				q			<=			16'h2C23;
		end
		32'h00008DD6: begin
				q			<=			16'h0001;
		end
		32'h00008DD8: begin
				q			<=			16'h0B93;
		end
		32'h00008DDA: begin
				q			<=			16'h0000;
		end
		32'h00008DDC: begin
				q			<=			16'h8413;
		end
		32'h00008DDE: begin
				q			<=			16'h0009;
		end
		32'h00008DE0: begin
				q			<=			16'h0693;
		end
		32'h00008DE2: begin
				q			<=			16'h0250;
		end
		32'h00008DE4: begin
				q			<=			16'h4783;
		end
		32'h00008DE6: begin
				q			<=			16'h0004;
		end
		32'h00008DE8: begin
				q			<=			16'h8463;
		end
		32'h00008DEA: begin
				q			<=			16'h0007;
		end
		32'h00008DEC: begin
				q			<=			16'h9663;
		end
		32'h00008DEE: begin
				q			<=			16'h0AD7;
		end
		32'h00008DF0: begin
				q			<=			16'h0A33;
		end
		32'h00008DF2: begin
				q			<=			16'h4134;
		end
		32'h00008DF4: begin
				q			<=			16'h0863;
		end
		32'h00008DF6: begin
				q			<=			16'h040A;
		end
		32'h00008DF8: begin
				q			<=			16'h2783;
		end
		32'h00008DFA: begin
				q			<=			16'h0481;
		end
		32'h00008DFC: begin
				q			<=			16'h2023;
		end
		32'h00008DFE: begin
				q			<=			16'h0137;
		end
		32'h00008E00: begin
				q			<=			16'h2223;
		end
		32'h00008E02: begin
				q			<=			16'h0147;
		end
		32'h00008E04: begin
				q			<=			16'h87B3;
		end
		32'h00008E06: begin
				q			<=			16'h0147;
		end
		32'h00008E08: begin
				q			<=			16'h2423;
		end
		32'h00008E0A: begin
				q			<=			16'h04F1;
		end
		32'h00008E0C: begin
				q			<=			16'h2783;
		end
		32'h00008E0E: begin
				q			<=			16'h0441;
		end
		32'h00008E10: begin
				q			<=			16'h0693;
		end
		32'h00008E12: begin
				q			<=			16'h0070;
		end
		32'h00008E14: begin
				q			<=			16'h0713;
		end
		32'h00008E16: begin
				q			<=			16'h0087;
		end
		32'h00008E18: begin
				q			<=			16'h8793;
		end
		32'h00008E1A: begin
				q			<=			16'h0017;
		end
		32'h00008E1C: begin
				q			<=			16'h2223;
		end
		32'h00008E1E: begin
				q			<=			16'h04F1;
		end
		32'h00008E20: begin
				q			<=			16'hD063;
		end
		32'h00008E22: begin
				q			<=			16'h02F6;
		end
		32'h00008E24: begin
				q			<=			16'h0613;
		end
		32'h00008E26: begin
				q			<=			16'h0401;
		end
		32'h00008E28: begin
				q			<=			16'h0593;
		end
		32'h00008E2A: begin
				q			<=			16'h0009;
		end
		32'h00008E2C: begin
				q			<=			16'h8513;
		end
		32'h00008E2E: begin
				q			<=			16'h000A;
		end
		32'h00008E30: begin
				q			<=			16'h0097;
		end
		32'h00008E32: begin
				q			<=			16'h0000;
		end
		32'h00008E34: begin
				q			<=			16'h80E7;
		end
		32'h00008E36: begin
				q			<=			16'hD2C0;
		end
		32'h00008E38: begin
				q			<=			16'h1CE3;
		end
		32'h00008E3A: begin
				q			<=			16'h2C05;
		end
		32'h00008E3C: begin
				q			<=			16'h0713;
		end
		32'h00008E3E: begin
				q			<=			16'h000B;
		end
		32'h00008E40: begin
				q			<=			16'h8BB3;
		end
		32'h00008E42: begin
				q			<=			16'h014B;
		end
		32'h00008E44: begin
				q			<=			16'h4783;
		end
		32'h00008E46: begin
				q			<=			16'h0004;
		end
		32'h00008E48: begin
				q			<=			16'h88E3;
		end
		32'h00008E4A: begin
				q			<=			16'h3407;
		end
		32'h00008E4C: begin
				q			<=			16'h0993;
		end
		32'h00008E4E: begin
				q			<=			16'h0014;
		end
		32'h00008E50: begin
				q			<=			16'h0DA3;
		end
		32'h00008E52: begin
				q			<=			16'h0201;
		end
		32'h00008E54: begin
				q			<=			16'h0413;
		end
		32'h00008E56: begin
				q			<=			16'hFFF0;
		end
		32'h00008E58: begin
				q			<=			16'h0A13;
		end
		32'h00008E5A: begin
				q			<=			16'h0000;
		end
		32'h00008E5C: begin
				q			<=			16'h0D13;
		end
		32'h00008E5E: begin
				q			<=			16'h0000;
		end
		32'h00008E60: begin
				q			<=			16'h0C13;
		end
		32'h00008E62: begin
				q			<=			16'h0090;
		end
		32'h00008E64: begin
				q			<=			16'h0513;
		end
		32'h00008E66: begin
				q			<=			16'h05A0;
		end
		32'h00008E68: begin
				q			<=			16'h0813;
		end
		32'h00008E6A: begin
				q			<=			16'h02A0;
		end
		32'h00008E6C: begin
				q			<=			16'hC603;
		end
		32'h00008E6E: begin
				q			<=			16'h0009;
		end
		32'h00008E70: begin
				q			<=			16'h8993;
		end
		32'h00008E72: begin
				q			<=			16'h0019;
		end
		32'h00008E74: begin
				q			<=			16'h0693;
		end
		32'h00008E76: begin
				q			<=			16'hFE06;
		end
		32'h00008E78: begin
				q			<=			16'h64E3;
		end
		32'h00008E7A: begin
				q			<=			16'h12D5;
		end
		32'h00008E7C: begin
				q			<=			16'h6797;
		end
		32'h00008E7E: begin
				q			<=			16'h0000;
		end
		32'h00008E80: begin
				q			<=			16'h8793;
		end
		32'h00008E82: begin
				q			<=			16'h7AC7;
		end
		32'h00008E84: begin
				q			<=			16'h9693;
		end
		32'h00008E86: begin
				q			<=			16'h0026;
		end
		32'h00008E88: begin
				q			<=			16'h86B3;
		end
		32'h00008E8A: begin
				q			<=			16'h00F6;
		end
		32'h00008E8C: begin
				q			<=			16'hA683;
		end
		32'h00008E8E: begin
				q			<=			16'h0006;
		end
		32'h00008E90: begin
				q			<=			16'h86B3;
		end
		32'h00008E92: begin
				q			<=			16'h00F6;
		end
		32'h00008E94: begin
				q			<=			16'h8067;
		end
		32'h00008E96: begin
				q			<=			16'h0006;
		end
		32'h00008E98: begin
				q			<=			16'h0413;
		end
		32'h00008E9A: begin
				q			<=			16'h0014;
		end
		32'h00008E9C: begin
				q			<=			16'hF06F;
		end
		32'h00008E9E: begin
				q			<=			16'hF49F;
		end
		32'h00008EA0: begin
				q			<=			16'h7797;
		end
		32'h00008EA2: begin
				q			<=			16'h0000;
		end
		32'h00008EA4: begin
				q			<=			16'h8793;
		end
		32'h00008EA6: begin
				q			<=			16'hEF87;
		end
		32'h00008EA8: begin
				q			<=			16'h2A23;
		end
		32'h00008EAA: begin
				q			<=			16'h00F1;
		end
		32'h00008EAC: begin
				q			<=			16'h7693;
		end
		32'h00008EAE: begin
				q			<=			16'h020D;
		end
		32'h00008EB0: begin
				q			<=			16'h8C63;
		end
		32'h00008EB2: begin
				q			<=			16'h6E06;
		end
		32'h00008EB4: begin
				q			<=			16'h8493;
		end
		32'h00008EB6: begin
				q			<=			16'h0074;
		end
		32'h00008EB8: begin
				q			<=			16'hF493;
		end
		32'h00008EBA: begin
				q			<=			16'hFF84;
		end
		32'h00008EBC: begin
				q			<=			16'hA883;
		end
		32'h00008EBE: begin
				q			<=			16'h0004;
		end
		32'h00008EC0: begin
				q			<=			16'hAC83;
		end
		32'h00008EC2: begin
				q			<=			16'h0044;
		end
		32'h00008EC4: begin
				q			<=			16'h8C13;
		end
		32'h00008EC6: begin
				q			<=			16'h0084;
		end
		32'h00008EC8: begin
				q			<=			16'h7693;
		end
		32'h00008ECA: begin
				q			<=			16'h001D;
		end
		32'h00008ECC: begin
				q			<=			16'h8E63;
		end
		32'h00008ECE: begin
				q			<=			16'h0006;
		end
		32'h00008ED0: begin
				q			<=			16'hE6B3;
		end
		32'h00008ED2: begin
				q			<=			16'h0198;
		end
		32'h00008ED4: begin
				q			<=			16'h8A63;
		end
		32'h00008ED6: begin
				q			<=			16'h0006;
		end
		32'h00008ED8: begin
				q			<=			16'h0693;
		end
		32'h00008EDA: begin
				q			<=			16'h0300;
		end
		32'h00008EDC: begin
				q			<=			16'h0E23;
		end
		32'h00008EDE: begin
				q			<=			16'h02D1;
		end
		32'h00008EE0: begin
				q			<=			16'h0EA3;
		end
		32'h00008EE2: begin
				q			<=			16'h02C1;
		end
		32'h00008EE4: begin
				q			<=			16'h6D13;
		end
		32'h00008EE6: begin
				q			<=			16'h002D;
		end
		32'h00008EE8: begin
				q			<=			16'h7D13;
		end
		32'h00008EEA: begin
				q			<=			16'hBFFD;
		end
		32'h00008EEC: begin
				q			<=			16'h006F;
		end
		32'h00008EEE: begin
				q			<=			16'h3280;
		end
		32'h00008EF0: begin
				q			<=			16'h8513;
		end
		32'h00008EF2: begin
				q			<=			16'h000A;
		end
		32'h00008EF4: begin
				q			<=			16'h2423;
		end
		32'h00008EF6: begin
				q			<=			16'h00E1;
		end
		32'h00008EF8: begin
				q			<=			16'hE0EF;
		end
		32'h00008EFA: begin
				q			<=			16'hC5CF;
		end
		32'h00008EFC: begin
				q			<=			16'h2783;
		end
		32'h00008EFE: begin
				q			<=			16'h0045;
		end
		32'h00008F00: begin
				q			<=			16'h8513;
		end
		32'h00008F02: begin
				q			<=			16'h0007;
		end
		32'h00008F04: begin
				q			<=			16'h2C23;
		end
		32'h00008F06: begin
				q			<=			16'h00F1;
		end
		32'h00008F08: begin
				q			<=			16'hA097;
		end
		32'h00008F0A: begin
				q			<=			16'hFFFF;
		end
		32'h00008F0C: begin
				q			<=			16'h80E7;
		end
		32'h00008F0E: begin
				q			<=			16'hF240;
		end
		32'h00008F10: begin
				q			<=			16'h2823;
		end
		32'h00008F12: begin
				q			<=			16'h00A1;
		end
		32'h00008F14: begin
				q			<=			16'h8513;
		end
		32'h00008F16: begin
				q			<=			16'h000A;
		end
		32'h00008F18: begin
				q			<=			16'hE0EF;
		end
		32'h00008F1A: begin
				q			<=			16'hC3CF;
		end
		32'h00008F1C: begin
				q			<=			16'h2783;
		end
		32'h00008F1E: begin
				q			<=			16'h0085;
		end
		32'h00008F20: begin
				q			<=			16'h2703;
		end
		32'h00008F22: begin
				q			<=			16'h0081;
		end
		32'h00008F24: begin
				q			<=			16'h2623;
		end
		32'h00008F26: begin
				q			<=			16'h00F1;
		end
		32'h00008F28: begin
				q			<=			16'h2783;
		end
		32'h00008F2A: begin
				q			<=			16'h0101;
		end
		32'h00008F2C: begin
				q			<=			16'h8CE3;
		end
		32'h00008F2E: begin
				q			<=			16'hF207;
		end
		32'h00008F30: begin
				q			<=			16'h2783;
		end
		32'h00008F32: begin
				q			<=			16'h00C1;
		end
		32'h00008F34: begin
				q			<=			16'h88E3;
		end
		32'h00008F36: begin
				q			<=			16'hF207;
		end
		32'h00008F38: begin
				q			<=			16'hC683;
		end
		32'h00008F3A: begin
				q			<=			16'h0007;
		end
		32'h00008F3C: begin
				q			<=			16'h84E3;
		end
		32'h00008F3E: begin
				q			<=			16'hF206;
		end
		32'h00008F40: begin
				q			<=			16'h6D13;
		end
		32'h00008F42: begin
				q			<=			16'h400D;
		end
		32'h00008F44: begin
				q			<=			16'hF06F;
		end
		32'h00008F46: begin
				q			<=			16'hF21F;
		end
		32'h00008F48: begin
				q			<=			16'h4683;
		end
		32'h00008F4A: begin
				q			<=			16'h03B1;
		end
		32'h00008F4C: begin
				q			<=			16'h9CE3;
		end
		32'h00008F4E: begin
				q			<=			16'hF006;
		end
		32'h00008F50: begin
				q			<=			16'h0693;
		end
		32'h00008F52: begin
				q			<=			16'h0200;
		end
		32'h00008F54: begin
				q			<=			16'h0DA3;
		end
		32'h00008F56: begin
				q			<=			16'h02D1;
		end
		32'h00008F58: begin
				q			<=			16'hF06F;
		end
		32'h00008F5A: begin
				q			<=			16'hF0DF;
		end
		32'h00008F5C: begin
				q			<=			16'h6D13;
		end
		32'h00008F5E: begin
				q			<=			16'h001D;
		end
		32'h00008F60: begin
				q			<=			16'hF06F;
		end
		32'h00008F62: begin
				q			<=			16'hF05F;
		end
		32'h00008F64: begin
				q			<=			16'hAA03;
		end
		32'h00008F66: begin
				q			<=			16'h0004;
		end
		32'h00008F68: begin
				q			<=			16'h8493;
		end
		32'h00008F6A: begin
				q			<=			16'h0044;
		end
		32'h00008F6C: begin
				q			<=			16'h5CE3;
		end
		32'h00008F6E: begin
				q			<=			16'hEE0A;
		end
		32'h00008F70: begin
				q			<=			16'h0A33;
		end
		32'h00008F72: begin
				q			<=			16'h4140;
		end
		32'h00008F74: begin
				q			<=			16'h6D13;
		end
		32'h00008F76: begin
				q			<=			16'h004D;
		end
		32'h00008F78: begin
				q			<=			16'hF06F;
		end
		32'h00008F7A: begin
				q			<=			16'hEEDF;
		end
		32'h00008F7C: begin
				q			<=			16'h0693;
		end
		32'h00008F7E: begin
				q			<=			16'h02B0;
		end
		32'h00008F80: begin
				q			<=			16'hF06F;
		end
		32'h00008F82: begin
				q			<=			16'hFD5F;
		end
		32'h00008F84: begin
				q			<=			16'hC603;
		end
		32'h00008F86: begin
				q			<=			16'h0009;
		end
		32'h00008F88: begin
				q			<=			16'h8693;
		end
		32'h00008F8A: begin
				q			<=			16'h0019;
		end
		32'h00008F8C: begin
				q			<=			16'h1263;
		end
		32'h00008F8E: begin
				q			<=			16'h0506;
		end
		32'h00008F90: begin
				q			<=			16'hA403;
		end
		32'h00008F92: begin
				q			<=			16'h0004;
		end
		32'h00008F94: begin
				q			<=			16'h8613;
		end
		32'h00008F96: begin
				q			<=			16'h0044;
		end
		32'h00008F98: begin
				q			<=			16'h5463;
		end
		32'h00008F9A: begin
				q			<=			16'h0004;
		end
		32'h00008F9C: begin
				q			<=			16'h0413;
		end
		32'h00008F9E: begin
				q			<=			16'hFFF0;
		end
		32'h00008FA0: begin
				q			<=			16'h0493;
		end
		32'h00008FA2: begin
				q			<=			16'h0006;
		end
		32'h00008FA4: begin
				q			<=			16'h8993;
		end
		32'h00008FA6: begin
				q			<=			16'h0006;
		end
		32'h00008FA8: begin
				q			<=			16'hF06F;
		end
		32'h00008FAA: begin
				q			<=			16'hEBDF;
		end
		32'h00008FAC: begin
				q			<=			16'h0793;
		end
		32'h00008FAE: begin
				q			<=			16'h00A0;
		end
		32'h00008FB0: begin
				q			<=			16'h0433;
		end
		32'h00008FB2: begin
				q			<=			16'h02F4;
		end
		32'h00008FB4: begin
				q			<=			16'h8693;
		end
		32'h00008FB6: begin
				q			<=			16'h0016;
		end
		32'h00008FB8: begin
				q			<=			16'hC603;
		end
		32'h00008FBA: begin
				q			<=			16'hFFF6;
		end
		32'h00008FBC: begin
				q			<=			16'h0433;
		end
		32'h00008FBE: begin
				q			<=			16'h00B4;
		end
		32'h00008FC0: begin
				q			<=			16'h0593;
		end
		32'h00008FC2: begin
				q			<=			16'hFD06;
		end
		32'h00008FC4: begin
				q			<=			16'h74E3;
		end
		32'h00008FC6: begin
				q			<=			16'hFEBC;
		end
		32'h00008FC8: begin
				q			<=			16'h8993;
		end
		32'h00008FCA: begin
				q			<=			16'h0006;
		end
		32'h00008FCC: begin
				q			<=			16'hF06F;
		end
		32'h00008FCE: begin
				q			<=			16'hEA9F;
		end
		32'h00008FD0: begin
				q			<=			16'h0413;
		end
		32'h00008FD2: begin
				q			<=			16'h0000;
		end
		32'h00008FD4: begin
				q			<=			16'hF06F;
		end
		32'h00008FD6: begin
				q			<=			16'hFEDF;
		end
		32'h00008FD8: begin
				q			<=			16'h6D13;
		end
		32'h00008FDA: begin
				q			<=			16'h080D;
		end
		32'h00008FDC: begin
				q			<=			16'hF06F;
		end
		32'h00008FDE: begin
				q			<=			16'hE89F;
		end
		32'h00008FE0: begin
				q			<=			16'h8693;
		end
		32'h00008FE2: begin
				q			<=			16'h0009;
		end
		32'h00008FE4: begin
				q			<=			16'h0A13;
		end
		32'h00008FE6: begin
				q			<=			16'h0000;
		end
		32'h00008FE8: begin
				q			<=			16'h0793;
		end
		32'h00008FEA: begin
				q			<=			16'h00A0;
		end
		32'h00008FEC: begin
				q			<=			16'h0A33;
		end
		32'h00008FEE: begin
				q			<=			16'h02FA;
		end
		32'h00008FF0: begin
				q			<=			16'h0613;
		end
		32'h00008FF2: begin
				q			<=			16'hFD06;
		end
		32'h00008FF4: begin
				q			<=			16'h8693;
		end
		32'h00008FF6: begin
				q			<=			16'h0016;
		end
		32'h00008FF8: begin
				q			<=			16'h0A33;
		end
		32'h00008FFA: begin
				q			<=			16'h0146;
		end
		32'h00008FFC: begin
				q			<=			16'hC603;
		end
		32'h00008FFE: begin
				q			<=			16'hFFF6;
		end
		32'h00009000: begin
				q			<=			16'h0593;
		end
		32'h00009002: begin
				q			<=			16'hFD06;
		end
		32'h00009004: begin
				q			<=			16'h72E3;
		end
		32'h00009006: begin
				q			<=			16'hFEBC;
		end
		32'h00009008: begin
				q			<=			16'hF06F;
		end
		32'h0000900A: begin
				q			<=			16'hFC1F;
		end
		32'h0000900C: begin
				q			<=			16'hC603;
		end
		32'h0000900E: begin
				q			<=			16'h0009;
		end
		32'h00009010: begin
				q			<=			16'h0693;
		end
		32'h00009012: begin
				q			<=			16'h0680;
		end
		32'h00009014: begin
				q			<=			16'h1863;
		end
		32'h00009016: begin
				q			<=			16'h00D6;
		end
		32'h00009018: begin
				q			<=			16'h8993;
		end
		32'h0000901A: begin
				q			<=			16'h0019;
		end
		32'h0000901C: begin
				q			<=			16'h6D13;
		end
		32'h0000901E: begin
				q			<=			16'h200D;
		end
		32'h00009020: begin
				q			<=			16'hF06F;
		end
		32'h00009022: begin
				q			<=			16'hE45F;
		end
		32'h00009024: begin
				q			<=			16'h6D13;
		end
		32'h00009026: begin
				q			<=			16'h040D;
		end
		32'h00009028: begin
				q			<=			16'hF06F;
		end
		32'h0000902A: begin
				q			<=			16'hE3DF;
		end
		32'h0000902C: begin
				q			<=			16'hC603;
		end
		32'h0000902E: begin
				q			<=			16'h0009;
		end
		32'h00009030: begin
				q			<=			16'h0693;
		end
		32'h00009032: begin
				q			<=			16'h06C0;
		end
		32'h00009034: begin
				q			<=			16'h1863;
		end
		32'h00009036: begin
				q			<=			16'h00D6;
		end
		32'h00009038: begin
				q			<=			16'h8993;
		end
		32'h0000903A: begin
				q			<=			16'h0019;
		end
		32'h0000903C: begin
				q			<=			16'h6D13;
		end
		32'h0000903E: begin
				q			<=			16'h020D;
		end
		32'h00009040: begin
				q			<=			16'hF06F;
		end
		32'h00009042: begin
				q			<=			16'hE25F;
		end
		32'h00009044: begin
				q			<=			16'h6D13;
		end
		32'h00009046: begin
				q			<=			16'h010D;
		end
		32'h00009048: begin
				q			<=			16'hF06F;
		end
		32'h0000904A: begin
				q			<=			16'hE1DF;
		end
		32'h0000904C: begin
				q			<=			16'hA683;
		end
		32'h0000904E: begin
				q			<=			16'h0004;
		end
		32'h00009050: begin
				q			<=			16'h8C13;
		end
		32'h00009052: begin
				q			<=			16'h0044;
		end
		32'h00009054: begin
				q			<=			16'h0DA3;
		end
		32'h00009056: begin
				q			<=			16'h0201;
		end
		32'h00009058: begin
				q			<=			16'h0623;
		end
		32'h0000905A: begin
				q			<=			16'h08D1;
		end
		32'h0000905C: begin
				q			<=			16'h0413;
		end
		32'h0000905E: begin
				q			<=			16'h0010;
		end
		32'h00009060: begin
				q			<=			16'h0C93;
		end
		32'h00009062: begin
				q			<=			16'h0000;
		end
		32'h00009064: begin
				q			<=			16'h0493;
		end
		32'h00009066: begin
				q			<=			16'h08C1;
		end
		32'h00009068: begin
				q			<=			16'h006F;
		end
		32'h0000906A: begin
				q			<=			16'h1F00;
		end
		32'h0000906C: begin
				q			<=			16'h6D13;
		end
		32'h0000906E: begin
				q			<=			16'h010D;
		end
		32'h00009070: begin
				q			<=			16'h7693;
		end
		32'h00009072: begin
				q			<=			16'h020D;
		end
		32'h00009074: begin
				q			<=			16'h8C63;
		end
		32'h00009076: begin
				q			<=			16'h0406;
		end
		32'h00009078: begin
				q			<=			16'h8493;
		end
		32'h0000907A: begin
				q			<=			16'h0074;
		end
		32'h0000907C: begin
				q			<=			16'hF493;
		end
		32'h0000907E: begin
				q			<=			16'hFF84;
		end
		32'h00009080: begin
				q			<=			16'hA883;
		end
		32'h00009082: begin
				q			<=			16'h0004;
		end
		32'h00009084: begin
				q			<=			16'hAC83;
		end
		32'h00009086: begin
				q			<=			16'h0044;
		end
		32'h00009088: begin
				q			<=			16'h8C13;
		end
		32'h0000908A: begin
				q			<=			16'h0084;
		end
		32'h0000908C: begin
				q			<=			16'hDE63;
		end
		32'h0000908E: begin
				q			<=			16'h000C;
		end
		32'h00009090: begin
				q			<=			16'h08B3;
		end
		32'h00009092: begin
				q			<=			16'h4110;
		end
		32'h00009094: begin
				q			<=			16'h36B3;
		end
		32'h00009096: begin
				q			<=			16'h0110;
		end
		32'h00009098: begin
				q			<=			16'h0333;
		end
		32'h0000909A: begin
				q			<=			16'h4190;
		end
		32'h0000909C: begin
				q			<=			16'h0CB3;
		end
		32'h0000909E: begin
				q			<=			16'h40D3;
		end
		32'h000090A0: begin
				q			<=			16'h0693;
		end
		32'h000090A2: begin
				q			<=			16'h02D0;
		end
		32'h000090A4: begin
				q			<=			16'h0DA3;
		end
		32'h000090A6: begin
				q			<=			16'h02D1;
		end
		32'h000090A8: begin
				q			<=			16'h0693;
		end
		32'h000090AA: begin
				q			<=			16'hFFF0;
		end
		32'h000090AC: begin
				q			<=			16'h1A63;
		end
		32'h000090AE: begin
				q			<=			16'h52D4;
		end
		32'h000090B0: begin
				q			<=			16'h9463;
		end
		32'h000090B2: begin
				q			<=			16'h5A0C;
		end
		32'h000090B4: begin
				q			<=			16'h0693;
		end
		32'h000090B6: begin
				q			<=			16'h0090;
		end
		32'h000090B8: begin
				q			<=			16'hE063;
		end
		32'h000090BA: begin
				q			<=			16'h5B16;
		end
		32'h000090BC: begin
				q			<=			16'h8893;
		end
		32'h000090BE: begin
				q			<=			16'h0308;
		end
		32'h000090C0: begin
				q			<=			16'h07A3;
		end
		32'h000090C2: begin
				q			<=			16'h0F11;
		end
		32'h000090C4: begin
				q			<=			16'h0493;
		end
		32'h000090C6: begin
				q			<=			16'h0EF1;
		end
		32'h000090C8: begin
				q			<=			16'h006F;
		end
		32'h000090CA: begin
				q			<=			16'h5780;
		end
		32'h000090CC: begin
				q			<=			16'h7693;
		end
		32'h000090CE: begin
				q			<=			16'h010D;
		end
		32'h000090D0: begin
				q			<=			16'h8C13;
		end
		32'h000090D2: begin
				q			<=			16'h0044;
		end
		32'h000090D4: begin
				q			<=			16'h8863;
		end
		32'h000090D6: begin
				q			<=			16'h0006;
		end
		32'h000090D8: begin
				q			<=			16'hA883;
		end
		32'h000090DA: begin
				q			<=			16'h0004;
		end
		32'h000090DC: begin
				q			<=			16'hDC93;
		end
		32'h000090DE: begin
				q			<=			16'h41F8;
		end
		32'h000090E0: begin
				q			<=			16'hF06F;
		end
		32'h000090E2: begin
				q			<=			16'hFADF;
		end
		32'h000090E4: begin
				q			<=			16'h7693;
		end
		32'h000090E6: begin
				q			<=			16'h040D;
		end
		32'h000090E8: begin
				q			<=			16'hA883;
		end
		32'h000090EA: begin
				q			<=			16'h0004;
		end
		32'h000090EC: begin
				q			<=			16'h8863;
		end
		32'h000090EE: begin
				q			<=			16'h0006;
		end
		32'h000090F0: begin
				q			<=			16'h9893;
		end
		32'h000090F2: begin
				q			<=			16'h0108;
		end
		32'h000090F4: begin
				q			<=			16'hD893;
		end
		32'h000090F6: begin
				q			<=			16'h4108;
		end
		32'h000090F8: begin
				q			<=			16'hF06F;
		end
		32'h000090FA: begin
				q			<=			16'hFE5F;
		end
		32'h000090FC: begin
				q			<=			16'h7693;
		end
		32'h000090FE: begin
				q			<=			16'h200D;
		end
		32'h00009100: begin
				q			<=			16'h8EE3;
		end
		32'h00009102: begin
				q			<=			16'hFC06;
		end
		32'h00009104: begin
				q			<=			16'h9893;
		end
		32'h00009106: begin
				q			<=			16'h0188;
		end
		32'h00009108: begin
				q			<=			16'hD893;
		end
		32'h0000910A: begin
				q			<=			16'h4188;
		end
		32'h0000910C: begin
				q			<=			16'hF06F;
		end
		32'h0000910E: begin
				q			<=			16'hFD1F;
		end
		32'h00009110: begin
				q			<=			16'h7613;
		end
		32'h00009112: begin
				q			<=			16'h020D;
		end
		32'h00009114: begin
				q			<=			16'hA683;
		end
		32'h00009116: begin
				q			<=			16'h0004;
		end
		32'h00009118: begin
				q			<=			16'h8493;
		end
		32'h0000911A: begin
				q			<=			16'h0044;
		end
		32'h0000911C: begin
				q			<=			16'h0A63;
		end
		32'h0000911E: begin
				q			<=			16'h0006;
		end
		32'h00009120: begin
				q			<=			16'hD793;
		end
		32'h00009122: begin
				q			<=			16'h41FB;
		end
		32'h00009124: begin
				q			<=			16'hA023;
		end
		32'h00009126: begin
				q			<=			16'h0176;
		end
		32'h00009128: begin
				q			<=			16'hA223;
		end
		32'h0000912A: begin
				q			<=			16'h00F6;
		end
		32'h0000912C: begin
				q			<=			16'hF06F;
		end
		32'h0000912E: begin
				q			<=			16'hCB1F;
		end
		32'h00009130: begin
				q			<=			16'h7613;
		end
		32'h00009132: begin
				q			<=			16'h010D;
		end
		32'h00009134: begin
				q			<=			16'h0663;
		end
		32'h00009136: begin
				q			<=			16'h0006;
		end
		32'h00009138: begin
				q			<=			16'hA023;
		end
		32'h0000913A: begin
				q			<=			16'h0176;
		end
		32'h0000913C: begin
				q			<=			16'hF06F;
		end
		32'h0000913E: begin
				q			<=			16'hCA1F;
		end
		32'h00009140: begin
				q			<=			16'h7613;
		end
		32'h00009142: begin
				q			<=			16'h040D;
		end
		32'h00009144: begin
				q			<=			16'h0663;
		end
		32'h00009146: begin
				q			<=			16'h0006;
		end
		32'h00009148: begin
				q			<=			16'h9023;
		end
		32'h0000914A: begin
				q			<=			16'h0176;
		end
		32'h0000914C: begin
				q			<=			16'hF06F;
		end
		32'h0000914E: begin
				q			<=			16'hC91F;
		end
		32'h00009150: begin
				q			<=			16'h7793;
		end
		32'h00009152: begin
				q			<=			16'h200D;
		end
		32'h00009154: begin
				q			<=			16'h82E3;
		end
		32'h00009156: begin
				q			<=			16'hFE07;
		end
		32'h00009158: begin
				q			<=			16'h8023;
		end
		32'h0000915A: begin
				q			<=			16'h0176;
		end
		32'h0000915C: begin
				q			<=			16'hF06F;
		end
		32'h0000915E: begin
				q			<=			16'hC81F;
		end
		32'h00009160: begin
				q			<=			16'h6D13;
		end
		32'h00009162: begin
				q			<=			16'h010D;
		end
		32'h00009164: begin
				q			<=			16'h7693;
		end
		32'h00009166: begin
				q			<=			16'h020D;
		end
		32'h00009168: begin
				q			<=			16'h8663;
		end
		32'h0000916A: begin
				q			<=			16'h0406;
		end
		32'h0000916C: begin
				q			<=			16'h8493;
		end
		32'h0000916E: begin
				q			<=			16'h0074;
		end
		32'h00009170: begin
				q			<=			16'hF493;
		end
		32'h00009172: begin
				q			<=			16'hFF84;
		end
		32'h00009174: begin
				q			<=			16'hA883;
		end
		32'h00009176: begin
				q			<=			16'h0004;
		end
		32'h00009178: begin
				q			<=			16'hAC83;
		end
		32'h0000917A: begin
				q			<=			16'h0044;
		end
		32'h0000917C: begin
				q			<=			16'h8C13;
		end
		32'h0000917E: begin
				q			<=			16'h0084;
		end
		32'h00009180: begin
				q			<=			16'h7D13;
		end
		32'h00009182: begin
				q			<=			16'hBFFD;
		end
		32'h00009184: begin
				q			<=			16'h0693;
		end
		32'h00009186: begin
				q			<=			16'h0000;
		end
		32'h00009188: begin
				q			<=			16'h0DA3;
		end
		32'h0000918A: begin
				q			<=			16'h0201;
		end
		32'h0000918C: begin
				q			<=			16'h0613;
		end
		32'h0000918E: begin
				q			<=			16'hFFF0;
		end
		32'h00009190: begin
				q			<=			16'h0E63;
		end
		32'h00009192: begin
				q			<=			16'h44C4;
		end
		32'h00009194: begin
				q			<=			16'h0613;
		end
		32'h00009196: begin
				q			<=			16'h000D;
		end
		32'h00009198: begin
				q			<=			16'hE5B3;
		end
		32'h0000919A: begin
				q			<=			16'h0198;
		end
		32'h0000919C: begin
				q			<=			16'h7D13;
		end
		32'h0000919E: begin
				q			<=			16'hF7FD;
		end
		32'h000091A0: begin
				q			<=			16'h9663;
		end
		32'h000091A2: begin
				q			<=			16'h4405;
		end
		32'h000091A4: begin
				q			<=			16'h0063;
		end
		32'h000091A6: begin
				q			<=			16'h5E04;
		end
		32'h000091A8: begin
				q			<=			16'h0613;
		end
		32'h000091AA: begin
				q			<=			16'h0010;
		end
		32'h000091AC: begin
				q			<=			16'h9463;
		end
		32'h000091AE: begin
				q			<=			16'h44C6;
		end
		32'h000091B0: begin
				q			<=			16'hF06F;
		end
		32'h000091B2: begin
				q			<=			16'hF0DF;
		end
		32'h000091B4: begin
				q			<=			16'h7693;
		end
		32'h000091B6: begin
				q			<=			16'h010D;
		end
		32'h000091B8: begin
				q			<=			16'h8C13;
		end
		32'h000091BA: begin
				q			<=			16'h0044;
		end
		32'h000091BC: begin
				q			<=			16'h8663;
		end
		32'h000091BE: begin
				q			<=			16'h0006;
		end
		32'h000091C0: begin
				q			<=			16'hA883;
		end
		32'h000091C2: begin
				q			<=			16'h0004;
		end
		32'h000091C4: begin
				q			<=			16'h006F;
		end
		32'h000091C6: begin
				q			<=			16'h0100;
		end
		32'h000091C8: begin
				q			<=			16'h7693;
		end
		32'h000091CA: begin
				q			<=			16'h040D;
		end
		32'h000091CC: begin
				q			<=			16'h8863;
		end
		32'h000091CE: begin
				q			<=			16'h0006;
		end
		32'h000091D0: begin
				q			<=			16'hD883;
		end
		32'h000091D2: begin
				q			<=			16'h0004;
		end
		32'h000091D4: begin
				q			<=			16'h0C93;
		end
		32'h000091D6: begin
				q			<=			16'h0000;
		end
		32'h000091D8: begin
				q			<=			16'hF06F;
		end
		32'h000091DA: begin
				q			<=			16'hFA9F;
		end
		32'h000091DC: begin
				q			<=			16'h7693;
		end
		32'h000091DE: begin
				q			<=			16'h200D;
		end
		32'h000091E0: begin
				q			<=			16'h80E3;
		end
		32'h000091E2: begin
				q			<=			16'hFE06;
		end
		32'h000091E4: begin
				q			<=			16'hC883;
		end
		32'h000091E6: begin
				q			<=			16'h0004;
		end
		32'h000091E8: begin
				q			<=			16'hF06F;
		end
		32'h000091EA: begin
				q			<=			16'hFEDF;
		end
		32'h000091EC: begin
				q			<=			16'h86B7;
		end
		32'h000091EE: begin
				q			<=			16'hFFFF;
		end
		32'h000091F0: begin
				q			<=			16'hA883;
		end
		32'h000091F2: begin
				q			<=			16'h0004;
		end
		32'h000091F4: begin
				q			<=			16'hC693;
		end
		32'h000091F6: begin
				q			<=			16'h8306;
		end
		32'h000091F8: begin
				q			<=			16'h7797;
		end
		32'h000091FA: begin
				q			<=			16'h0000;
		end
		32'h000091FC: begin
				q			<=			16'h8793;
		end
		32'h000091FE: begin
				q			<=			16'hB8C7;
		end
		32'h00009200: begin
				q			<=			16'h8C13;
		end
		32'h00009202: begin
				q			<=			16'h0044;
		end
		32'h00009204: begin
				q			<=			16'h0C93;
		end
		32'h00009206: begin
				q			<=			16'h0000;
		end
		32'h00009208: begin
				q			<=			16'h6D13;
		end
		32'h0000920A: begin
				q			<=			16'h002D;
		end
		32'h0000920C: begin
				q			<=			16'h1E23;
		end
		32'h0000920E: begin
				q			<=			16'h02D1;
		end
		32'h00009210: begin
				q			<=			16'h2A23;
		end
		32'h00009212: begin
				q			<=			16'h00F1;
		end
		32'h00009214: begin
				q			<=			16'h0693;
		end
		32'h00009216: begin
				q			<=			16'h0020;
		end
		32'h00009218: begin
				q			<=			16'hF06F;
		end
		32'h0000921A: begin
				q			<=			16'hF71F;
		end
		32'h0000921C: begin
				q			<=			16'h0DA3;
		end
		32'h0000921E: begin
				q			<=			16'h0201;
		end
		32'h00009220: begin
				q			<=			16'h0693;
		end
		32'h00009222: begin
				q			<=			16'hFFF0;
		end
		32'h00009224: begin
				q			<=			16'h2423;
		end
		32'h00009226: begin
				q			<=			16'h00E1;
		end
		32'h00009228: begin
				q			<=			16'h8C13;
		end
		32'h0000922A: begin
				q			<=			16'h0044;
		end
		32'h0000922C: begin
				q			<=			16'hA483;
		end
		32'h0000922E: begin
				q			<=			16'h0004;
		end
		32'h00009230: begin
				q			<=			16'h0863;
		end
		32'h00009232: begin
				q			<=			16'h2ED4;
		end
		32'h00009234: begin
				q			<=			16'h0613;
		end
		32'h00009236: begin
				q			<=			16'h0004;
		end
		32'h00009238: begin
				q			<=			16'h0593;
		end
		32'h0000923A: begin
				q			<=			16'h0000;
		end
		32'h0000923C: begin
				q			<=			16'h8513;
		end
		32'h0000923E: begin
				q			<=			16'h0004;
		end
		32'h00009240: begin
				q			<=			16'hF097;
		end
		32'h00009242: begin
				q			<=			16'hFFFF;
		end
		32'h00009244: begin
				q			<=			16'h80E7;
		end
		32'h00009246: begin
				q			<=			16'h8180;
		end
		32'h00009248: begin
				q			<=			16'h0C93;
		end
		32'h0000924A: begin
				q			<=			16'h0000;
		end
		32'h0000924C: begin
				q			<=			16'h2703;
		end
		32'h0000924E: begin
				q			<=			16'h0081;
		end
		32'h00009250: begin
				q			<=			16'h0463;
		end
		32'h00009252: begin
				q			<=			16'h0005;
		end
		32'h00009254: begin
				q			<=			16'h0433;
		end
		32'h00009256: begin
				q			<=			16'h4095;
		end
		32'h00009258: begin
				q			<=			16'h2423;
		end
		32'h0000925A: begin
				q			<=			16'h0191;
		end
		32'h0000925C: begin
				q			<=			16'hD463;
		end
		32'h0000925E: begin
				q			<=			16'h008C;
		end
		32'h00009260: begin
				q			<=			16'h2423;
		end
		32'h00009262: begin
				q			<=			16'h0081;
		end
		32'h00009264: begin
				q			<=			16'h4683;
		end
		32'h00009266: begin
				q			<=			16'h03B1;
		end
		32'h00009268: begin
				q			<=			16'h8863;
		end
		32'h0000926A: begin
				q			<=			16'h0006;
		end
		32'h0000926C: begin
				q			<=			16'h2783;
		end
		32'h0000926E: begin
				q			<=			16'h0081;
		end
		32'h00009270: begin
				q			<=			16'h8793;
		end
		32'h00009272: begin
				q			<=			16'h0017;
		end
		32'h00009274: begin
				q			<=			16'h2423;
		end
		32'h00009276: begin
				q			<=			16'h00F1;
		end
		32'h00009278: begin
				q			<=			16'h7D93;
		end
		32'h0000927A: begin
				q			<=			16'h002D;
		end
		32'h0000927C: begin
				q			<=			16'h8863;
		end
		32'h0000927E: begin
				q			<=			16'h000D;
		end
		32'h00009280: begin
				q			<=			16'h2783;
		end
		32'h00009282: begin
				q			<=			16'h0081;
		end
		32'h00009284: begin
				q			<=			16'h8793;
		end
		32'h00009286: begin
				q			<=			16'h0027;
		end
		32'h00009288: begin
				q			<=			16'h2423;
		end
		32'h0000928A: begin
				q			<=			16'h00F1;
		end
		32'h0000928C: begin
				q			<=			16'h7793;
		end
		32'h0000928E: begin
				q			<=			16'h084D;
		end
		32'h00009290: begin
				q			<=			16'h2E23;
		end
		32'h00009292: begin
				q			<=			16'h00F1;
		end
		32'h00009294: begin
				q			<=			16'h9863;
		end
		32'h00009296: begin
				q			<=			16'h0607;
		end
		32'h00009298: begin
				q			<=			16'h2783;
		end
		32'h0000929A: begin
				q			<=			16'h0081;
		end
		32'h0000929C: begin
				q			<=			16'h06B3;
		end
		32'h0000929E: begin
				q			<=			16'h40FA;
		end
		32'h000092A0: begin
				q			<=			16'h5263;
		end
		32'h000092A2: begin
				q			<=			16'h06D0;
		end
		32'h000092A4: begin
				q			<=			16'h0893;
		end
		32'h000092A6: begin
				q			<=			16'h0100;
		end
		32'h000092A8: begin
				q			<=			16'h6817;
		end
		32'h000092AA: begin
				q			<=			16'h0000;
		end
		32'h000092AC: begin
				q			<=			16'h0813;
		end
		32'h000092AE: begin
				q			<=			16'h4EC8;
		end
		32'h000092B0: begin
				q			<=			16'h0313;
		end
		32'h000092B2: begin
				q			<=			16'h0070;
		end
		32'h000092B4: begin
				q			<=			16'h2603;
		end
		32'h000092B6: begin
				q			<=			16'h0441;
		end
		32'h000092B8: begin
				q			<=			16'h2023;
		end
		32'h000092BA: begin
				q			<=			16'h0107;
		end
		32'h000092BC: begin
				q			<=			16'h2583;
		end
		32'h000092BE: begin
				q			<=			16'h0481;
		end
		32'h000092C0: begin
				q			<=			16'h0613;
		end
		32'h000092C2: begin
				q			<=			16'h0016;
		end
		32'h000092C4: begin
				q			<=			16'h0513;
		end
		32'h000092C6: begin
				q			<=			16'h0087;
		end
		32'h000092C8: begin
				q			<=			16'hC663;
		end
		32'h000092CA: begin
				q			<=			16'h4ED8;
		end
		32'h000092CC: begin
				q			<=			16'h2223;
		end
		32'h000092CE: begin
				q			<=			16'h00D7;
		end
		32'h000092D0: begin
				q			<=			16'h86B3;
		end
		32'h000092D2: begin
				q			<=			16'h00B6;
		end
		32'h000092D4: begin
				q			<=			16'h2423;
		end
		32'h000092D6: begin
				q			<=			16'h04D1;
		end
		32'h000092D8: begin
				q			<=			16'h2223;
		end
		32'h000092DA: begin
				q			<=			16'h04C1;
		end
		32'h000092DC: begin
				q			<=			16'h0693;
		end
		32'h000092DE: begin
				q			<=			16'h0070;
		end
		32'h000092E0: begin
				q			<=			16'h0713;
		end
		32'h000092E2: begin
				q			<=			16'h0005;
		end
		32'h000092E4: begin
				q			<=			16'hD063;
		end
		32'h000092E6: begin
				q			<=			16'h02C6;
		end
		32'h000092E8: begin
				q			<=			16'h0613;
		end
		32'h000092EA: begin
				q			<=			16'h0401;
		end
		32'h000092EC: begin
				q			<=			16'h0593;
		end
		32'h000092EE: begin
				q			<=			16'h0009;
		end
		32'h000092F0: begin
				q			<=			16'h8513;
		end
		32'h000092F2: begin
				q			<=			16'h000A;
		end
		32'h000092F4: begin
				q			<=			16'h0097;
		end
		32'h000092F6: begin
				q			<=			16'h0000;
		end
		32'h000092F8: begin
				q			<=			16'h80E7;
		end
		32'h000092FA: begin
				q			<=			16'h8680;
		end
		32'h000092FC: begin
				q			<=			16'h1A63;
		end
		32'h000092FE: begin
				q			<=			16'h6005;
		end
		32'h00009300: begin
				q			<=			16'h0713;
		end
		32'h00009302: begin
				q			<=			16'h000B;
		end
		32'h00009304: begin
				q			<=			16'h4683;
		end
		32'h00009306: begin
				q			<=			16'h03B1;
		end
		32'h00009308: begin
				q			<=			16'h8A63;
		end
		32'h0000930A: begin
				q			<=			16'h0406;
		end
		32'h0000930C: begin
				q			<=			16'h0613;
		end
		32'h0000930E: begin
				q			<=			16'h03B1;
		end
		32'h00009310: begin
				q			<=			16'h2023;
		end
		32'h00009312: begin
				q			<=			16'h00C7;
		end
		32'h00009314: begin
				q			<=			16'h0613;
		end
		32'h00009316: begin
				q			<=			16'h0010;
		end
		32'h00009318: begin
				q			<=			16'h2683;
		end
		32'h0000931A: begin
				q			<=			16'h0441;
		end
		32'h0000931C: begin
				q			<=			16'h2223;
		end
		32'h0000931E: begin
				q			<=			16'h00C7;
		end
		32'h00009320: begin
				q			<=			16'h2603;
		end
		32'h00009322: begin
				q			<=			16'h0481;
		end
		32'h00009324: begin
				q			<=			16'h8693;
		end
		32'h00009326: begin
				q			<=			16'h0016;
		end
		32'h00009328: begin
				q			<=			16'h2223;
		end
		32'h0000932A: begin
				q			<=			16'h04D1;
		end
		32'h0000932C: begin
				q			<=			16'h0613;
		end
		32'h0000932E: begin
				q			<=			16'h0016;
		end
		32'h00009330: begin
				q			<=			16'h2423;
		end
		32'h00009332: begin
				q			<=			16'h04C1;
		end
		32'h00009334: begin
				q			<=			16'h0613;
		end
		32'h00009336: begin
				q			<=			16'h0070;
		end
		32'h00009338: begin
				q			<=			16'h0713;
		end
		32'h0000933A: begin
				q			<=			16'h0087;
		end
		32'h0000933C: begin
				q			<=			16'h5063;
		end
		32'h0000933E: begin
				q			<=			16'h02D6;
		end
		32'h00009340: begin
				q			<=			16'h0613;
		end
		32'h00009342: begin
				q			<=			16'h0401;
		end
		32'h00009344: begin
				q			<=			16'h0593;
		end
		32'h00009346: begin
				q			<=			16'h0009;
		end
		32'h00009348: begin
				q			<=			16'h8513;
		end
		32'h0000934A: begin
				q			<=			16'h000A;
		end
		32'h0000934C: begin
				q			<=			16'h0097;
		end
		32'h0000934E: begin
				q			<=			16'h0000;
		end
		32'h00009350: begin
				q			<=			16'h80E7;
		end
		32'h00009352: begin
				q			<=			16'h8100;
		end
		32'h00009354: begin
				q			<=			16'h1E63;
		end
		32'h00009356: begin
				q			<=			16'h5A05;
		end
		32'h00009358: begin
				q			<=			16'h0713;
		end
		32'h0000935A: begin
				q			<=			16'h000B;
		end
		32'h0000935C: begin
				q			<=			16'h8A63;
		end
		32'h0000935E: begin
				q			<=			16'h040D;
		end
		32'h00009360: begin
				q			<=			16'h0613;
		end
		32'h00009362: begin
				q			<=			16'h03C1;
		end
		32'h00009364: begin
				q			<=			16'h2023;
		end
		32'h00009366: begin
				q			<=			16'h00C7;
		end
		32'h00009368: begin
				q			<=			16'h0613;
		end
		32'h0000936A: begin
				q			<=			16'h0020;
		end
		32'h0000936C: begin
				q			<=			16'h2683;
		end
		32'h0000936E: begin
				q			<=			16'h0441;
		end
		32'h00009370: begin
				q			<=			16'h2223;
		end
		32'h00009372: begin
				q			<=			16'h00C7;
		end
		32'h00009374: begin
				q			<=			16'h2603;
		end
		32'h00009376: begin
				q			<=			16'h0481;
		end
		32'h00009378: begin
				q			<=			16'h8693;
		end
		32'h0000937A: begin
				q			<=			16'h0016;
		end
		32'h0000937C: begin
				q			<=			16'h2223;
		end
		32'h0000937E: begin
				q			<=			16'h04D1;
		end
		32'h00009380: begin
				q			<=			16'h0613;
		end
		32'h00009382: begin
				q			<=			16'h0026;
		end
		32'h00009384: begin
				q			<=			16'h2423;
		end
		32'h00009386: begin
				q			<=			16'h04C1;
		end
		32'h00009388: begin
				q			<=			16'h0613;
		end
		32'h0000938A: begin
				q			<=			16'h0070;
		end
		32'h0000938C: begin
				q			<=			16'h0713;
		end
		32'h0000938E: begin
				q			<=			16'h0087;
		end
		32'h00009390: begin
				q			<=			16'h5063;
		end
		32'h00009392: begin
				q			<=			16'h02D6;
		end
		32'h00009394: begin
				q			<=			16'h0613;
		end
		32'h00009396: begin
				q			<=			16'h0401;
		end
		32'h00009398: begin
				q			<=			16'h0593;
		end
		32'h0000939A: begin
				q			<=			16'h0009;
		end
		32'h0000939C: begin
				q			<=			16'h8513;
		end
		32'h0000939E: begin
				q			<=			16'h000A;
		end
		32'h000093A0: begin
				q			<=			16'hF097;
		end
		32'h000093A2: begin
				q			<=			16'hFFFF;
		end
		32'h000093A4: begin
				q			<=			16'h80E7;
		end
		32'h000093A6: begin
				q			<=			16'h7BC0;
		end
		32'h000093A8: begin
				q			<=			16'h1463;
		end
		32'h000093AA: begin
				q			<=			16'h5605;
		end
		32'h000093AC: begin
				q			<=			16'h0713;
		end
		32'h000093AE: begin
				q			<=			16'h000B;
		end
		32'h000093B0: begin
				q			<=			16'h2783;
		end
		32'h000093B2: begin
				q			<=			16'h01C1;
		end
		32'h000093B4: begin
				q			<=			16'h0693;
		end
		32'h000093B6: begin
				q			<=			16'h0800;
		end
		32'h000093B8: begin
				q			<=			16'h9863;
		end
		32'h000093BA: begin
				q			<=			16'h06D7;
		end
		32'h000093BC: begin
				q			<=			16'h2783;
		end
		32'h000093BE: begin
				q			<=			16'h0081;
		end
		32'h000093C0: begin
				q			<=			16'h0DB3;
		end
		32'h000093C2: begin
				q			<=			16'h40FA;
		end
		32'h000093C4: begin
				q			<=			16'h5263;
		end
		32'h000093C6: begin
				q			<=			16'h07B0;
		end
		32'h000093C8: begin
				q			<=			16'h0893;
		end
		32'h000093CA: begin
				q			<=			16'h0100;
		end
		32'h000093CC: begin
				q			<=			16'h6817;
		end
		32'h000093CE: begin
				q			<=			16'h0000;
		end
		32'h000093D0: begin
				q			<=			16'h0813;
		end
		32'h000093D2: begin
				q			<=			16'h3D88;
		end
		32'h000093D4: begin
				q			<=			16'h0313;
		end
		32'h000093D6: begin
				q			<=			16'h0070;
		end
		32'h000093D8: begin
				q			<=			16'h2683;
		end
		32'h000093DA: begin
				q			<=			16'h0441;
		end
		32'h000093DC: begin
				q			<=			16'h2023;
		end
		32'h000093DE: begin
				q			<=			16'h0107;
		end
		32'h000093E0: begin
				q			<=			16'h2603;
		end
		32'h000093E2: begin
				q			<=			16'h0481;
		end
		32'h000093E4: begin
				q			<=			16'h8693;
		end
		32'h000093E6: begin
				q			<=			16'h0016;
		end
		32'h000093E8: begin
				q			<=			16'h0593;
		end
		32'h000093EA: begin
				q			<=			16'h0087;
		end
		32'h000093EC: begin
				q			<=			16'hC263;
		end
		32'h000093EE: begin
				q			<=			16'h43B8;
		end
		32'h000093F0: begin
				q			<=			16'h0633;
		end
		32'h000093F2: begin
				q			<=			16'h01B6;
		end
		32'h000093F4: begin
				q			<=			16'h2223;
		end
		32'h000093F6: begin
				q			<=			16'h01B7;
		end
		32'h000093F8: begin
				q			<=			16'h2423;
		end
		32'h000093FA: begin
				q			<=			16'h04C1;
		end
		32'h000093FC: begin
				q			<=			16'h2223;
		end
		32'h000093FE: begin
				q			<=			16'h04D1;
		end
		32'h00009400: begin
				q			<=			16'h0613;
		end
		32'h00009402: begin
				q			<=			16'h0070;
		end
		32'h00009404: begin
				q			<=			16'h8713;
		end
		32'h00009406: begin
				q			<=			16'h0005;
		end
		32'h00009408: begin
				q			<=			16'h5063;
		end
		32'h0000940A: begin
				q			<=			16'h02D6;
		end
		32'h0000940C: begin
				q			<=			16'h0613;
		end
		32'h0000940E: begin
				q			<=			16'h0401;
		end
		32'h00009410: begin
				q			<=			16'h0593;
		end
		32'h00009412: begin
				q			<=			16'h0009;
		end
		32'h00009414: begin
				q			<=			16'h8513;
		end
		32'h00009416: begin
				q			<=			16'h000A;
		end
		32'h00009418: begin
				q			<=			16'hF097;
		end
		32'h0000941A: begin
				q			<=			16'hFFFF;
		end
		32'h0000941C: begin
				q			<=			16'h80E7;
		end
		32'h0000941E: begin
				q			<=			16'h7440;
		end
		32'h00009420: begin
				q			<=			16'h1863;
		end
		32'h00009422: begin
				q			<=			16'h4E05;
		end
		32'h00009424: begin
				q			<=			16'h0713;
		end
		32'h00009426: begin
				q			<=			16'h000B;
		end
		32'h00009428: begin
				q			<=			16'h8CB3;
		end
		32'h0000942A: begin
				q			<=			16'h408C;
		end
		32'h0000942C: begin
				q			<=			16'h5263;
		end
		32'h0000942E: begin
				q			<=			16'h0790;
		end
		32'h00009430: begin
				q			<=			16'h0813;
		end
		32'h00009432: begin
				q			<=			16'h0100;
		end
		32'h00009434: begin
				q			<=			16'h6D97;
		end
		32'h00009436: begin
				q			<=			16'h0000;
		end
		32'h00009438: begin
				q			<=			16'h8D93;
		end
		32'h0000943A: begin
				q			<=			16'h370D;
		end
		32'h0000943C: begin
				q			<=			16'h0893;
		end
		32'h0000943E: begin
				q			<=			16'h0070;
		end
		32'h00009440: begin
				q			<=			16'h2683;
		end
		32'h00009442: begin
				q			<=			16'h0441;
		end
		32'h00009444: begin
				q			<=			16'h2023;
		end
		32'h00009446: begin
				q			<=			16'h01B7;
		end
		32'h00009448: begin
				q			<=			16'h2603;
		end
		32'h0000944A: begin
				q			<=			16'h0481;
		end
		32'h0000944C: begin
				q			<=			16'h8693;
		end
		32'h0000944E: begin
				q			<=			16'h0016;
		end
		32'h00009450: begin
				q			<=			16'h0593;
		end
		32'h00009452: begin
				q			<=			16'h0087;
		end
		32'h00009454: begin
				q			<=			16'h4863;
		end
		32'h00009456: begin
				q			<=			16'h4198;
		end
		32'h00009458: begin
				q			<=			16'h2223;
		end
		32'h0000945A: begin
				q			<=			16'h0197;
		end
		32'h0000945C: begin
				q			<=			16'h8CB3;
		end
		32'h0000945E: begin
				q			<=			16'h00CC;
		end
		32'h00009460: begin
				q			<=			16'h2423;
		end
		32'h00009462: begin
				q			<=			16'h0591;
		end
		32'h00009464: begin
				q			<=			16'h2223;
		end
		32'h00009466: begin
				q			<=			16'h04D1;
		end
		32'h00009468: begin
				q			<=			16'h0613;
		end
		32'h0000946A: begin
				q			<=			16'h0070;
		end
		32'h0000946C: begin
				q			<=			16'h8713;
		end
		32'h0000946E: begin
				q			<=			16'h0005;
		end
		32'h00009470: begin
				q			<=			16'h5063;
		end
		32'h00009472: begin
				q			<=			16'h02D6;
		end
		32'h00009474: begin
				q			<=			16'h0613;
		end
		32'h00009476: begin
				q			<=			16'h0401;
		end
		32'h00009478: begin
				q			<=			16'h0593;
		end
		32'h0000947A: begin
				q			<=			16'h0009;
		end
		32'h0000947C: begin
				q			<=			16'h8513;
		end
		32'h0000947E: begin
				q			<=			16'h000A;
		end
		32'h00009480: begin
				q			<=			16'hF097;
		end
		32'h00009482: begin
				q			<=			16'hFFFF;
		end
		32'h00009484: begin
				q			<=			16'h80E7;
		end
		32'h00009486: begin
				q			<=			16'h6DC0;
		end
		32'h00009488: begin
				q			<=			16'h1463;
		end
		32'h0000948A: begin
				q			<=			16'h4805;
		end
		32'h0000948C: begin
				q			<=			16'h0713;
		end
		32'h0000948E: begin
				q			<=			16'h000B;
		end
		32'h00009490: begin
				q			<=			16'h2683;
		end
		32'h00009492: begin
				q			<=			16'h0481;
		end
		32'h00009494: begin
				q			<=			16'h2223;
		end
		32'h00009496: begin
				q			<=			16'h0087;
		end
		32'h00009498: begin
				q			<=			16'h2023;
		end
		32'h0000949A: begin
				q			<=			16'h0097;
		end
		32'h0000949C: begin
				q			<=			16'h8433;
		end
		32'h0000949E: begin
				q			<=			16'h0086;
		end
		32'h000094A0: begin
				q			<=			16'h2683;
		end
		32'h000094A2: begin
				q			<=			16'h0441;
		end
		32'h000094A4: begin
				q			<=			16'h2423;
		end
		32'h000094A6: begin
				q			<=			16'h0481;
		end
		32'h000094A8: begin
				q			<=			16'h0613;
		end
		32'h000094AA: begin
				q			<=			16'h0070;
		end
		32'h000094AC: begin
				q			<=			16'h8693;
		end
		32'h000094AE: begin
				q			<=			16'h0016;
		end
		32'h000094B0: begin
				q			<=			16'h2223;
		end
		32'h000094B2: begin
				q			<=			16'h04D1;
		end
		32'h000094B4: begin
				q			<=			16'h0713;
		end
		32'h000094B6: begin
				q			<=			16'h0087;
		end
		32'h000094B8: begin
				q			<=			16'h5063;
		end
		32'h000094BA: begin
				q			<=			16'h02D6;
		end
		32'h000094BC: begin
				q			<=			16'h0613;
		end
		32'h000094BE: begin
				q			<=			16'h0401;
		end
		32'h000094C0: begin
				q			<=			16'h0593;
		end
		32'h000094C2: begin
				q			<=			16'h0009;
		end
		32'h000094C4: begin
				q			<=			16'h8513;
		end
		32'h000094C6: begin
				q			<=			16'h000A;
		end
		32'h000094C8: begin
				q			<=			16'hF097;
		end
		32'h000094CA: begin
				q			<=			16'hFFFF;
		end
		32'h000094CC: begin
				q			<=			16'h80E7;
		end
		32'h000094CE: begin
				q			<=			16'h6940;
		end
		32'h000094D0: begin
				q			<=			16'h1063;
		end
		32'h000094D2: begin
				q			<=			16'h4405;
		end
		32'h000094D4: begin
				q			<=			16'h0713;
		end
		32'h000094D6: begin
				q			<=			16'h000B;
		end
		32'h000094D8: begin
				q			<=			16'h7793;
		end
		32'h000094DA: begin
				q			<=			16'h004D;
		end
		32'h000094DC: begin
				q			<=			16'h9A63;
		end
		32'h000094DE: begin
				q			<=			16'h3C07;
		end
		32'h000094E0: begin
				q			<=			16'h2783;
		end
		32'h000094E2: begin
				q			<=			16'h0081;
		end
		32'h000094E4: begin
				q			<=			16'h5463;
		end
		32'h000094E6: begin
				q			<=			16'h00FA;
		end
		32'h000094E8: begin
				q			<=			16'h8A13;
		end
		32'h000094EA: begin
				q			<=			16'h0007;
		end
		32'h000094EC: begin
				q			<=			16'h2783;
		end
		32'h000094EE: begin
				q			<=			16'h0481;
		end
		32'h000094F0: begin
				q			<=			16'h8BB3;
		end
		32'h000094F2: begin
				q			<=			16'h014B;
		end
		32'h000094F4: begin
				q			<=			16'h8E63;
		end
		32'h000094F6: begin
				q			<=			16'h0007;
		end
		32'h000094F8: begin
				q			<=			16'h0613;
		end
		32'h000094FA: begin
				q			<=			16'h0401;
		end
		32'h000094FC: begin
				q			<=			16'h0593;
		end
		32'h000094FE: begin
				q			<=			16'h0009;
		end
		32'h00009500: begin
				q			<=			16'h8513;
		end
		32'h00009502: begin
				q			<=			16'h000A;
		end
		32'h00009504: begin
				q			<=			16'hF097;
		end
		32'h00009506: begin
				q			<=			16'hFFFF;
		end
		32'h00009508: begin
				q			<=			16'h80E7;
		end
		32'h0000950A: begin
				q			<=			16'h6580;
		end
		32'h0000950C: begin
				q			<=			16'h1263;
		end
		32'h0000950E: begin
				q			<=			16'h4005;
		end
		32'h00009510: begin
				q			<=			16'h2223;
		end
		32'h00009512: begin
				q			<=			16'h0401;
		end
		32'h00009514: begin
				q			<=			16'h0493;
		end
		32'h00009516: begin
				q			<=			16'h000C;
		end
		32'h00009518: begin
				q			<=			16'h0713;
		end
		32'h0000951A: begin
				q			<=			16'h000B;
		end
		32'h0000951C: begin
				q			<=			16'hF06F;
		end
		32'h0000951E: begin
				q			<=			16'h8C1F;
		end
		32'h00009520: begin
				q			<=			16'h8513;
		end
		32'h00009522: begin
				q			<=			16'h0004;
		end
		32'h00009524: begin
				q			<=			16'hA097;
		end
		32'h00009526: begin
				q			<=			16'hFFFF;
		end
		32'h00009528: begin
				q			<=			16'h80E7;
		end
		32'h0000952A: begin
				q			<=			16'h9080;
		end
		32'h0000952C: begin
				q			<=			16'h0413;
		end
		32'h0000952E: begin
				q			<=			16'h0005;
		end
		32'h00009530: begin
				q			<=			16'h0C93;
		end
		32'h00009532: begin
				q			<=			16'h0000;
		end
		32'h00009534: begin
				q			<=			16'h2703;
		end
		32'h00009536: begin
				q			<=			16'h0081;
		end
		32'h00009538: begin
				q			<=			16'hF06F;
		end
		32'h0000953A: begin
				q			<=			16'hD21F;
		end
		32'h0000953C: begin
				q			<=			16'h6D13;
		end
		32'h0000953E: begin
				q			<=			16'h010D;
		end
		32'h00009540: begin
				q			<=			16'h7693;
		end
		32'h00009542: begin
				q			<=			16'h020D;
		end
		32'h00009544: begin
				q			<=			16'h8063;
		end
		32'h00009546: begin
				q			<=			16'h0206;
		end
		32'h00009548: begin
				q			<=			16'h8493;
		end
		32'h0000954A: begin
				q			<=			16'h0074;
		end
		32'h0000954C: begin
				q			<=			16'hF493;
		end
		32'h0000954E: begin
				q			<=			16'hFF84;
		end
		32'h00009550: begin
				q			<=			16'hA883;
		end
		32'h00009552: begin
				q			<=			16'h0004;
		end
		32'h00009554: begin
				q			<=			16'hAC83;
		end
		32'h00009556: begin
				q			<=			16'h0044;
		end
		32'h00009558: begin
				q			<=			16'h8C13;
		end
		32'h0000955A: begin
				q			<=			16'h0084;
		end
		32'h0000955C: begin
				q			<=			16'h0693;
		end
		32'h0000955E: begin
				q			<=			16'h0010;
		end
		32'h00009560: begin
				q			<=			16'hF06F;
		end
		32'h00009562: begin
				q			<=			16'hC29F;
		end
		32'h00009564: begin
				q			<=			16'h7693;
		end
		32'h00009566: begin
				q			<=			16'h010D;
		end
		32'h00009568: begin
				q			<=			16'h8C13;
		end
		32'h0000956A: begin
				q			<=			16'h0044;
		end
		32'h0000956C: begin
				q			<=			16'h8663;
		end
		32'h0000956E: begin
				q			<=			16'h0006;
		end
		32'h00009570: begin
				q			<=			16'hA883;
		end
		32'h00009572: begin
				q			<=			16'h0004;
		end
		32'h00009574: begin
				q			<=			16'h006F;
		end
		32'h00009576: begin
				q			<=			16'h0100;
		end
		32'h00009578: begin
				q			<=			16'h7693;
		end
		32'h0000957A: begin
				q			<=			16'h040D;
		end
		32'h0000957C: begin
				q			<=			16'h8863;
		end
		32'h0000957E: begin
				q			<=			16'h0006;
		end
		32'h00009580: begin
				q			<=			16'hD883;
		end
		32'h00009582: begin
				q			<=			16'h0004;
		end
		32'h00009584: begin
				q			<=			16'h0C93;
		end
		32'h00009586: begin
				q			<=			16'h0000;
		end
		32'h00009588: begin
				q			<=			16'hF06F;
		end
		32'h0000958A: begin
				q			<=			16'hFD5F;
		end
		32'h0000958C: begin
				q			<=			16'h7693;
		end
		32'h0000958E: begin
				q			<=			16'h200D;
		end
		32'h00009590: begin
				q			<=			16'h80E3;
		end
		32'h00009592: begin
				q			<=			16'hFE06;
		end
		32'h00009594: begin
				q			<=			16'hC883;
		end
		32'h00009596: begin
				q			<=			16'h0004;
		end
		32'h00009598: begin
				q			<=			16'hF06F;
		end
		32'h0000959A: begin
				q			<=			16'hFEDF;
		end
		32'h0000959C: begin
				q			<=			16'h6797;
		end
		32'h0000959E: begin
				q			<=			16'h0000;
		end
		32'h000095A0: begin
				q			<=			16'h8793;
		end
		32'h000095A2: begin
				q			<=			16'h7E87;
		end
		32'h000095A4: begin
				q			<=			16'hF06F;
		end
		32'h000095A6: begin
				q			<=			16'h905F;
		end
		32'h000095A8: begin
				q			<=			16'h7693;
		end
		32'h000095AA: begin
				q			<=			16'h010D;
		end
		32'h000095AC: begin
				q			<=			16'h8C13;
		end
		32'h000095AE: begin
				q			<=			16'h0044;
		end
		32'h000095B0: begin
				q			<=			16'h8663;
		end
		32'h000095B2: begin
				q			<=			16'h0006;
		end
		32'h000095B4: begin
				q			<=			16'hA883;
		end
		32'h000095B6: begin
				q			<=			16'h0004;
		end
		32'h000095B8: begin
				q			<=			16'h006F;
		end
		32'h000095BA: begin
				q			<=			16'h0100;
		end
		32'h000095BC: begin
				q			<=			16'h7693;
		end
		32'h000095BE: begin
				q			<=			16'h040D;
		end
		32'h000095C0: begin
				q			<=			16'h8863;
		end
		32'h000095C2: begin
				q			<=			16'h0006;
		end
		32'h000095C4: begin
				q			<=			16'hD883;
		end
		32'h000095C6: begin
				q			<=			16'h0004;
		end
		32'h000095C8: begin
				q			<=			16'h0C93;
		end
		32'h000095CA: begin
				q			<=			16'h0000;
		end
		32'h000095CC: begin
				q			<=			16'hF06F;
		end
		32'h000095CE: begin
				q			<=			16'h8FDF;
		end
		32'h000095D0: begin
				q			<=			16'h7693;
		end
		32'h000095D2: begin
				q			<=			16'h200D;
		end
		32'h000095D4: begin
				q			<=			16'h80E3;
		end
		32'h000095D6: begin
				q			<=			16'hFE06;
		end
		32'h000095D8: begin
				q			<=			16'hC883;
		end
		32'h000095DA: begin
				q			<=			16'h0004;
		end
		32'h000095DC: begin
				q			<=			16'hF06F;
		end
		32'h000095DE: begin
				q			<=			16'hFEDF;
		end
		32'h000095E0: begin
				q			<=			16'h0613;
		end
		32'h000095E2: begin
				q			<=			16'h000D;
		end
		32'h000095E4: begin
				q			<=			16'h0693;
		end
		32'h000095E6: begin
				q			<=			16'h0010;
		end
		32'h000095E8: begin
				q			<=			16'hF06F;
		end
		32'h000095EA: begin
				q			<=			16'hBB1F;
		end
		32'h000095EC: begin
				q			<=			16'h0613;
		end
		32'h000095EE: begin
				q			<=			16'h0010;
		end
		32'h000095F0: begin
				q			<=			16'h80E3;
		end
		32'h000095F2: begin
				q			<=			16'hACC6;
		end
		32'h000095F4: begin
				q			<=			16'h0613;
		end
		32'h000095F6: begin
				q			<=			16'h0020;
		end
		32'h000095F8: begin
				q			<=			16'h8A63;
		end
		32'h000095FA: begin
				q			<=			16'h14C6;
		end
		32'h000095FC: begin
				q			<=			16'h0693;
		end
		32'h000095FE: begin
				q			<=			16'h0F01;
		end
		32'h00009600: begin
				q			<=			16'h9593;
		end
		32'h00009602: begin
				q			<=			16'h01DC;
		end
		32'h00009604: begin
				q			<=			16'hF613;
		end
		32'h00009606: begin
				q			<=			16'h0078;
		end
		32'h00009608: begin
				q			<=			16'hD893;
		end
		32'h0000960A: begin
				q			<=			16'h0038;
		end
		32'h0000960C: begin
				q			<=			16'h0613;
		end
		32'h0000960E: begin
				q			<=			16'h0306;
		end
		32'h00009610: begin
				q			<=			16'hE8B3;
		end
		32'h00009612: begin
				q			<=			16'h0115;
		end
		32'h00009614: begin
				q			<=			16'hDC93;
		end
		32'h00009616: begin
				q			<=			16'h003C;
		end
		32'h00009618: begin
				q			<=			16'h8FA3;
		end
		32'h0000961A: begin
				q			<=			16'hFEC6;
		end
		32'h0000961C: begin
				q			<=			16'hE5B3;
		end
		32'h0000961E: begin
				q			<=			16'h0198;
		end
		32'h00009620: begin
				q			<=			16'h8493;
		end
		32'h00009622: begin
				q			<=			16'hFFF6;
		end
		32'h00009624: begin
				q			<=			16'h9663;
		end
		32'h00009626: begin
				q			<=			16'h0205;
		end
		32'h00009628: begin
				q			<=			16'h7593;
		end
		32'h0000962A: begin
				q			<=			16'h001D;
		end
		32'h0000962C: begin
				q			<=			16'h8A63;
		end
		32'h0000962E: begin
				q			<=			16'h0005;
		end
		32'h00009630: begin
				q			<=			16'h0593;
		end
		32'h00009632: begin
				q			<=			16'h0300;
		end
		32'h00009634: begin
				q			<=			16'h0663;
		end
		32'h00009636: begin
				q			<=			16'h00B6;
		end
		32'h00009638: begin
				q			<=			16'h8FA3;
		end
		32'h0000963A: begin
				q			<=			16'hFEB4;
		end
		32'h0000963C: begin
				q			<=			16'h8493;
		end
		32'h0000963E: begin
				q			<=			16'hFFE6;
		end
		32'h00009640: begin
				q			<=			16'h0793;
		end
		32'h00009642: begin
				q			<=			16'h0F01;
		end
		32'h00009644: begin
				q			<=			16'h0C93;
		end
		32'h00009646: begin
				q			<=			16'h0004;
		end
		32'h00009648: begin
				q			<=			16'h8433;
		end
		32'h0000964A: begin
				q			<=			16'h4097;
		end
		32'h0000964C: begin
				q			<=			16'hF06F;
		end
		32'h0000964E: begin
				q			<=			16'hC0DF;
		end
		32'h00009650: begin
				q			<=			16'h8693;
		end
		32'h00009652: begin
				q			<=			16'h0004;
		end
		32'h00009654: begin
				q			<=			16'hF06F;
		end
		32'h00009656: begin
				q			<=			16'hFADF;
		end
		32'h00009658: begin
				q			<=			16'h7793;
		end
		32'h0000965A: begin
				q			<=			16'h400D;
		end
		32'h0000965C: begin
				q			<=			16'h0D93;
		end
		32'h0000965E: begin
				q			<=			16'h0000;
		end
		32'h00009660: begin
				q			<=			16'h0E13;
		end
		32'h00009662: begin
				q			<=			16'h0F01;
		end
		32'h00009664: begin
				q			<=			16'h2423;
		end
		32'h00009666: begin
				q			<=			16'h00F1;
		end
		32'h00009668: begin
				q			<=			16'h8513;
		end
		32'h0000966A: begin
				q			<=			16'h0008;
		end
		32'h0000966C: begin
				q			<=			16'h0613;
		end
		32'h0000966E: begin
				q			<=			16'h00A0;
		end
		32'h00009670: begin
				q			<=			16'h0693;
		end
		32'h00009672: begin
				q			<=			16'h0000;
		end
		32'h00009674: begin
				q			<=			16'h8593;
		end
		32'h00009676: begin
				q			<=			16'h000C;
		end
		32'h00009678: begin
				q			<=			16'h2223;
		end
		32'h0000967A: begin
				q			<=			16'h02E1;
		end
		32'h0000967C: begin
				q			<=			16'h0493;
		end
		32'h0000967E: begin
				q			<=			16'hFFFE;
		end
		32'h00009680: begin
				q			<=			16'h2023;
		end
		32'h00009682: begin
				q			<=			16'h03C1;
		end
		32'h00009684: begin
				q			<=			16'h2E23;
		end
		32'h00009686: begin
				q			<=			16'h0111;
		end
		32'h00009688: begin
				q			<=			16'h2097;
		end
		32'h0000968A: begin
				q			<=			16'h0000;
		end
		32'h0000968C: begin
				q			<=			16'h80E7;
		end
		32'h0000968E: begin
				q			<=			16'h85C0;
		end
		32'h00009690: begin
				q			<=			16'h2E03;
		end
		32'h00009692: begin
				q			<=			16'h0201;
		end
		32'h00009694: begin
				q			<=			16'h2783;
		end
		32'h00009696: begin
				q			<=			16'h0081;
		end
		32'h00009698: begin
				q			<=			16'h0513;
		end
		32'h0000969A: begin
				q			<=			16'h0305;
		end
		32'h0000969C: begin
				q			<=			16'h0FA3;
		end
		32'h0000969E: begin
				q			<=			16'hFEAE;
		end
		32'h000096A0: begin
				q			<=			16'h8D93;
		end
		32'h000096A2: begin
				q			<=			16'h001D;
		end
		32'h000096A4: begin
				q			<=			16'h2883;
		end
		32'h000096A6: begin
				q			<=			16'h01C1;
		end
		32'h000096A8: begin
				q			<=			16'h2703;
		end
		32'h000096AA: begin
				q			<=			16'h0241;
		end
		32'h000096AC: begin
				q			<=			16'h8463;
		end
		32'h000096AE: begin
				q			<=			16'h0607;
		end
		32'h000096B0: begin
				q			<=			16'h2783;
		end
		32'h000096B2: begin
				q			<=			16'h00C1;
		end
		32'h000096B4: begin
				q			<=			16'hC683;
		end
		32'h000096B6: begin
				q			<=			16'h0007;
		end
		32'h000096B8: begin
				q			<=			16'h9E63;
		end
		32'h000096BA: begin
				q			<=			16'h05B6;
		end
		32'h000096BC: begin
				q			<=			16'h0793;
		end
		32'h000096BE: begin
				q			<=			16'h0FF0;
		end
		32'h000096C0: begin
				q			<=			16'h8A63;
		end
		32'h000096C2: begin
				q			<=			16'h04FD;
		end
		32'h000096C4: begin
				q			<=			16'h9663;
		end
		32'h000096C6: begin
				q			<=			16'h000C;
		end
		32'h000096C8: begin
				q			<=			16'h0793;
		end
		32'h000096CA: begin
				q			<=			16'h0090;
		end
		32'h000096CC: begin
				q			<=			16'hF463;
		end
		32'h000096CE: begin
				q			<=			16'h0517;
		end
		32'h000096D0: begin
				q			<=			16'h2783;
		end
		32'h000096D2: begin
				q			<=			16'h0101;
		end
		32'h000096D4: begin
				q			<=			16'h2583;
		end
		32'h000096D6: begin
				q			<=			16'h0181;
		end
		32'h000096D8: begin
				q			<=			16'h2023;
		end
		32'h000096DA: begin
				q			<=			16'h0311;
		end
		32'h000096DC: begin
				q			<=			16'h84B3;
		end
		32'h000096DE: begin
				q			<=			16'h40F4;
		end
		32'h000096E0: begin
				q			<=			16'h8613;
		end
		32'h000096E2: begin
				q			<=			16'h0007;
		end
		32'h000096E4: begin
				q			<=			16'h8513;
		end
		32'h000096E6: begin
				q			<=			16'h0004;
		end
		32'h000096E8: begin
				q			<=			16'h2E23;
		end
		32'h000096EA: begin
				q			<=			16'h00E1;
		end
		32'h000096EC: begin
				q			<=			16'h9097;
		end
		32'h000096EE: begin
				q			<=			16'hFFFF;
		end
		32'h000096F0: begin
				q			<=			16'h80E7;
		end
		32'h000096F2: begin
				q			<=			16'h7A00;
		end
		32'h000096F4: begin
				q			<=			16'h2783;
		end
		32'h000096F6: begin
				q			<=			16'h00C1;
		end
		32'h000096F8: begin
				q			<=			16'h0D93;
		end
		32'h000096FA: begin
				q			<=			16'h0000;
		end
		32'h000096FC: begin
				q			<=			16'h2703;
		end
		32'h000096FE: begin
				q			<=			16'h01C1;
		end
		32'h00009700: begin
				q			<=			16'hC683;
		end
		32'h00009702: begin
				q			<=			16'h0017;
		end
		32'h00009704: begin
				q			<=			16'h2883;
		end
		32'h00009706: begin
				q			<=			16'h0201;
		end
		32'h00009708: begin
				q			<=			16'h8663;
		end
		32'h0000970A: begin
				q			<=			16'h0006;
		end
		32'h0000970C: begin
				q			<=			16'h8793;
		end
		32'h0000970E: begin
				q			<=			16'h0017;
		end
		32'h00009710: begin
				q			<=			16'h2623;
		end
		32'h00009712: begin
				q			<=			16'h00F1;
		end
		32'h00009714: begin
				q			<=			16'h8513;
		end
		32'h00009716: begin
				q			<=			16'h0008;
		end
		32'h00009718: begin
				q			<=			16'h8593;
		end
		32'h0000971A: begin
				q			<=			16'h000C;
		end
		32'h0000971C: begin
				q			<=			16'h0613;
		end
		32'h0000971E: begin
				q			<=			16'h00A0;
		end
		32'h00009720: begin
				q			<=			16'h0693;
		end
		32'h00009722: begin
				q			<=			16'h0000;
		end
		32'h00009724: begin
				q			<=			16'h2E23;
		end
		32'h00009726: begin
				q			<=			16'h00E1;
		end
		32'h00009728: begin
				q			<=			16'h1097;
		end
		32'h0000972A: begin
				q			<=			16'h0000;
		end
		32'h0000972C: begin
				q			<=			16'h80E7;
		end
		32'h0000972E: begin
				q			<=			16'h3840;
		end
		32'h00009730: begin
				q			<=			16'h8C93;
		end
		32'h00009732: begin
				q			<=			16'h0005;
		end
		32'h00009734: begin
				q			<=			16'hE5B3;
		end
		32'h00009736: begin
				q			<=			16'h00A5;
		end
		32'h00009738: begin
				q			<=			16'h0893;
		end
		32'h0000973A: begin
				q			<=			16'h0005;
		end
		32'h0000973C: begin
				q			<=			16'h2703;
		end
		32'h0000973E: begin
				q			<=			16'h01C1;
		end
		32'h00009740: begin
				q			<=			16'h80E3;
		end
		32'h00009742: begin
				q			<=			16'hF005;
		end
		32'h00009744: begin
				q			<=			16'h8E13;
		end
		32'h00009746: begin
				q			<=			16'h0004;
		end
		32'h00009748: begin
				q			<=			16'hF06F;
		end
		32'h0000974A: begin
				q			<=			16'hF21F;
		end
		32'h0000974C: begin
				q			<=			16'h0493;
		end
		32'h0000974E: begin
				q			<=			16'h0F01;
		end
		32'h00009750: begin
				q			<=			16'h2783;
		end
		32'h00009752: begin
				q			<=			16'h0141;
		end
		32'h00009754: begin
				q			<=			16'hF693;
		end
		32'h00009756: begin
				q			<=			16'h00F8;
		end
		32'h00009758: begin
				q			<=			16'h8493;
		end
		32'h0000975A: begin
				q			<=			16'hFFF4;
		end
		32'h0000975C: begin
				q			<=			16'h86B3;
		end
		32'h0000975E: begin
				q			<=			16'h00D7;
		end
		32'h00009760: begin
				q			<=			16'hC683;
		end
		32'h00009762: begin
				q			<=			16'h0006;
		end
		32'h00009764: begin
				q			<=			16'hD893;
		end
		32'h00009766: begin
				q			<=			16'h0048;
		end
		32'h00009768: begin
				q			<=			16'h8023;
		end
		32'h0000976A: begin
				q			<=			16'h00D4;
		end
		32'h0000976C: begin
				q			<=			16'h9693;
		end
		32'h0000976E: begin
				q			<=			16'h01CC;
		end
		32'h00009770: begin
				q			<=			16'hE8B3;
		end
		32'h00009772: begin
				q			<=			16'h0116;
		end
		32'h00009774: begin
				q			<=			16'hDC93;
		end
		32'h00009776: begin
				q			<=			16'h004C;
		end
		32'h00009778: begin
				q			<=			16'hE6B3;
		end
		32'h0000977A: begin
				q			<=			16'h0198;
		end
		32'h0000977C: begin
				q			<=			16'h9AE3;
		end
		32'h0000977E: begin
				q			<=			16'hFC06;
		end
		32'h00009780: begin
				q			<=			16'hF06F;
		end
		32'h00009782: begin
				q			<=			16'hEC1F;
		end
		32'h00009784: begin
				q			<=			16'h0493;
		end
		32'h00009786: begin
				q			<=			16'h0F01;
		end
		32'h00009788: begin
				q			<=			16'h9CE3;
		end
		32'h0000978A: begin
				q			<=			16'hEA06;
		end
		32'h0000978C: begin
				q			<=			16'h7613;
		end
		32'h0000978E: begin
				q			<=			16'h0016;
		end
		32'h00009790: begin
				q			<=			16'h08E3;
		end
		32'h00009792: begin
				q			<=			16'hEA06;
		end
		32'h00009794: begin
				q			<=			16'h0693;
		end
		32'h00009796: begin
				q			<=			16'h0300;
		end
		32'h00009798: begin
				q			<=			16'h07A3;
		end
		32'h0000979A: begin
				q			<=			16'h0ED1;
		end
		32'h0000979C: begin
				q			<=			16'hF06F;
		end
		32'h0000979E: begin
				q			<=			16'h929F;
		end
		32'h000097A0: begin
				q			<=			16'h0C63;
		end
		32'h000097A2: begin
				q			<=			16'h1E06;
		end
		32'h000097A4: begin
				q			<=			16'h0623;
		end
		32'h000097A6: begin
				q			<=			16'h08C1;
		end
		32'h000097A8: begin
				q			<=			16'h0DA3;
		end
		32'h000097AA: begin
				q			<=			16'h0201;
		end
		32'h000097AC: begin
				q			<=			16'h8C13;
		end
		32'h000097AE: begin
				q			<=			16'h0004;
		end
		32'h000097B0: begin
				q			<=			16'hF06F;
		end
		32'h000097B2: begin
				q			<=			16'h8ADF;
		end
		32'h000097B4: begin
				q			<=			16'h8593;
		end
		32'h000097B6: begin
				q			<=			16'h0105;
		end
		32'h000097B8: begin
				q			<=			16'h2223;
		end
		32'h000097BA: begin
				q			<=			16'h0117;
		end
		32'h000097BC: begin
				q			<=			16'h2423;
		end
		32'h000097BE: begin
				q			<=			16'h04B1;
		end
		32'h000097C0: begin
				q			<=			16'h2223;
		end
		32'h000097C2: begin
				q			<=			16'h04C1;
		end
		32'h000097C4: begin
				q			<=			16'h5063;
		end
		32'h000097C6: begin
				q			<=			16'h04C3;
		end
		32'h000097C8: begin
				q			<=			16'h0613;
		end
		32'h000097CA: begin
				q			<=			16'h0401;
		end
		32'h000097CC: begin
				q			<=			16'h0593;
		end
		32'h000097CE: begin
				q			<=			16'h0009;
		end
		32'h000097D0: begin
				q			<=			16'h8513;
		end
		32'h000097D2: begin
				q			<=			16'h000A;
		end
		32'h000097D4: begin
				q			<=			16'h2623;
		end
		32'h000097D6: begin
				q			<=			16'h0261;
		end
		32'h000097D8: begin
				q			<=			16'h2423;
		end
		32'h000097DA: begin
				q			<=			16'h0301;
		end
		32'h000097DC: begin
				q			<=			16'h2223;
		end
		32'h000097DE: begin
				q			<=			16'h0311;
		end
		32'h000097E0: begin
				q			<=			16'h2023;
		end
		32'h000097E2: begin
				q			<=			16'h02D1;
		end
		32'h000097E4: begin
				q			<=			16'hF097;
		end
		32'h000097E6: begin
				q			<=			16'hFFFF;
		end
		32'h000097E8: begin
				q			<=			16'h80E7;
		end
		32'h000097EA: begin
				q			<=			16'h3780;
		end
		32'h000097EC: begin
				q			<=			16'h1263;
		end
		32'h000097EE: begin
				q			<=			16'h1205;
		end
		32'h000097F0: begin
				q			<=			16'h2303;
		end
		32'h000097F2: begin
				q			<=			16'h02C1;
		end
		32'h000097F4: begin
				q			<=			16'h2803;
		end
		32'h000097F6: begin
				q			<=			16'h0281;
		end
		32'h000097F8: begin
				q			<=			16'h2883;
		end
		32'h000097FA: begin
				q			<=			16'h0241;
		end
		32'h000097FC: begin
				q			<=			16'h2683;
		end
		32'h000097FE: begin
				q			<=			16'h0201;
		end
		32'h00009800: begin
				q			<=			16'h0513;
		end
		32'h00009802: begin
				q			<=			16'h000B;
		end
		32'h00009804: begin
				q			<=			16'h8693;
		end
		32'h00009806: begin
				q			<=			16'hFF06;
		end
		32'h00009808: begin
				q			<=			16'h0713;
		end
		32'h0000980A: begin
				q			<=			16'h0005;
		end
		32'h0000980C: begin
				q			<=			16'hF06F;
		end
		32'h0000980E: begin
				q			<=			16'hAA9F;
		end
		32'h00009810: begin
				q			<=			16'h0613;
		end
		32'h00009812: begin
				q			<=			16'h0106;
		end
		32'h00009814: begin
				q			<=			16'h2223;
		end
		32'h00009816: begin
				q			<=			16'h0117;
		end
		32'h00009818: begin
				q			<=			16'h2423;
		end
		32'h0000981A: begin
				q			<=			16'h04C1;
		end
		32'h0000981C: begin
				q			<=			16'h2223;
		end
		32'h0000981E: begin
				q			<=			16'h04D1;
		end
		32'h00009820: begin
				q			<=			16'h5C63;
		end
		32'h00009822: begin
				q			<=			16'h02D3;
		end
		32'h00009824: begin
				q			<=			16'h0613;
		end
		32'h00009826: begin
				q			<=			16'h0401;
		end
		32'h00009828: begin
				q			<=			16'h0593;
		end
		32'h0000982A: begin
				q			<=			16'h0009;
		end
		32'h0000982C: begin
				q			<=			16'h8513;
		end
		32'h0000982E: begin
				q			<=			16'h000A;
		end
		32'h00009830: begin
				q			<=			16'h2223;
		end
		32'h00009832: begin
				q			<=			16'h0261;
		end
		32'h00009834: begin
				q			<=			16'h2023;
		end
		32'h00009836: begin
				q			<=			16'h0301;
		end
		32'h00009838: begin
				q			<=			16'h2E23;
		end
		32'h0000983A: begin
				q			<=			16'h0111;
		end
		32'h0000983C: begin
				q			<=			16'hF097;
		end
		32'h0000983E: begin
				q			<=			16'hFFFF;
		end
		32'h00009840: begin
				q			<=			16'h80E7;
		end
		32'h00009842: begin
				q			<=			16'h3200;
		end
		32'h00009844: begin
				q			<=			16'h1663;
		end
		32'h00009846: begin
				q			<=			16'h0C05;
		end
		32'h00009848: begin
				q			<=			16'h2303;
		end
		32'h0000984A: begin
				q			<=			16'h0241;
		end
		32'h0000984C: begin
				q			<=			16'h2803;
		end
		32'h0000984E: begin
				q			<=			16'h0201;
		end
		32'h00009850: begin
				q			<=			16'h2883;
		end
		32'h00009852: begin
				q			<=			16'h01C1;
		end
		32'h00009854: begin
				q			<=			16'h0593;
		end
		32'h00009856: begin
				q			<=			16'h000B;
		end
		32'h00009858: begin
				q			<=			16'h8D93;
		end
		32'h0000985A: begin
				q			<=			16'hFF0D;
		end
		32'h0000985C: begin
				q			<=			16'h8713;
		end
		32'h0000985E: begin
				q			<=			16'h0005;
		end
		32'h00009860: begin
				q			<=			16'hF06F;
		end
		32'h00009862: begin
				q			<=			16'hB79F;
		end
		32'h00009864: begin
				q			<=			16'h0613;
		end
		32'h00009866: begin
				q			<=			16'h0106;
		end
		32'h00009868: begin
				q			<=			16'h2223;
		end
		32'h0000986A: begin
				q			<=			16'h0107;
		end
		32'h0000986C: begin
				q			<=			16'h2423;
		end
		32'h0000986E: begin
				q			<=			16'h04C1;
		end
		32'h00009870: begin
				q			<=			16'h2223;
		end
		32'h00009872: begin
				q			<=			16'h04D1;
		end
		32'h00009874: begin
				q			<=			16'hD863;
		end
		32'h00009876: begin
				q			<=			16'h02D8;
		end
		32'h00009878: begin
				q			<=			16'h0613;
		end
		32'h0000987A: begin
				q			<=			16'h0401;
		end
		32'h0000987C: begin
				q			<=			16'h0593;
		end
		32'h0000987E: begin
				q			<=			16'h0009;
		end
		32'h00009880: begin
				q			<=			16'h8513;
		end
		32'h00009882: begin
				q			<=			16'h000A;
		end
		32'h00009884: begin
				q			<=			16'h2023;
		end
		32'h00009886: begin
				q			<=			16'h0311;
		end
		32'h00009888: begin
				q			<=			16'h2E23;
		end
		32'h0000988A: begin
				q			<=			16'h0101;
		end
		32'h0000988C: begin
				q			<=			16'hF097;
		end
		32'h0000988E: begin
				q			<=			16'hFFFF;
		end
		32'h00009890: begin
				q			<=			16'h80E7;
		end
		32'h00009892: begin
				q			<=			16'h2D00;
		end
		32'h00009894: begin
				q			<=			16'h1E63;
		end
		32'h00009896: begin
				q			<=			16'h0605;
		end
		32'h00009898: begin
				q			<=			16'h2883;
		end
		32'h0000989A: begin
				q			<=			16'h0201;
		end
		32'h0000989C: begin
				q			<=			16'h2803;
		end
		32'h0000989E: begin
				q			<=			16'h01C1;
		end
		32'h000098A0: begin
				q			<=			16'h0593;
		end
		32'h000098A2: begin
				q			<=			16'h000B;
		end
		32'h000098A4: begin
				q			<=			16'h8C93;
		end
		32'h000098A6: begin
				q			<=			16'hFF0C;
		end
		32'h000098A8: begin
				q			<=			16'h8713;
		end
		32'h000098AA: begin
				q			<=			16'h0005;
		end
		32'h000098AC: begin
				q			<=			16'hF06F;
		end
		32'h000098AE: begin
				q			<=			16'hB95F;
		end
		32'h000098B0: begin
				q			<=			16'h2783;
		end
		32'h000098B2: begin
				q			<=			16'h0081;
		end
		32'h000098B4: begin
				q			<=			16'h0433;
		end
		32'h000098B6: begin
				q			<=			16'h40FA;
		end
		32'h000098B8: begin
				q			<=			16'h54E3;
		end
		32'h000098BA: begin
				q			<=			16'hC280;
		end
		32'h000098BC: begin
				q			<=			16'h0C93;
		end
		32'h000098BE: begin
				q			<=			16'h0100;
		end
		32'h000098C0: begin
				q			<=			16'h6497;
		end
		32'h000098C2: begin
				q			<=			16'h0000;
		end
		32'h000098C4: begin
				q			<=			16'h8493;
		end
		32'h000098C6: begin
				q			<=			16'hED44;
		end
		32'h000098C8: begin
				q			<=			16'h0D93;
		end
		32'h000098CA: begin
				q			<=			16'h0070;
		end
		32'h000098CC: begin
				q			<=			16'h2783;
		end
		32'h000098CE: begin
				q			<=			16'h0441;
		end
		32'h000098D0: begin
				q			<=			16'h2023;
		end
		32'h000098D2: begin
				q			<=			16'h0097;
		end
		32'h000098D4: begin
				q			<=			16'h2683;
		end
		32'h000098D6: begin
				q			<=			16'h0481;
		end
		32'h000098D8: begin
				q			<=			16'h8793;
		end
		32'h000098DA: begin
				q			<=			16'h0017;
		end
		32'h000098DC: begin
				q			<=			16'hC063;
		end
		32'h000098DE: begin
				q			<=			16'h088C;
		end
		32'h000098E0: begin
				q			<=			16'h2223;
		end
		32'h000098E2: begin
				q			<=			16'h0087;
		end
		32'h000098E4: begin
				q			<=			16'h0433;
		end
		32'h000098E6: begin
				q			<=			16'h00D4;
		end
		32'h000098E8: begin
				q			<=			16'h2423;
		end
		32'h000098EA: begin
				q			<=			16'h0481;
		end
		32'h000098EC: begin
				q			<=			16'h2223;
		end
		32'h000098EE: begin
				q			<=			16'h04F1;
		end
		32'h000098F0: begin
				q			<=			16'h0713;
		end
		32'h000098F2: begin
				q			<=			16'h0070;
		end
		32'h000098F4: begin
				q			<=			16'h56E3;
		end
		32'h000098F6: begin
				q			<=			16'hBEF7;
		end
		32'h000098F8: begin
				q			<=			16'h0613;
		end
		32'h000098FA: begin
				q			<=			16'h0401;
		end
		32'h000098FC: begin
				q			<=			16'h0593;
		end
		32'h000098FE: begin
				q			<=			16'h0009;
		end
		32'h00009900: begin
				q			<=			16'h8513;
		end
		32'h00009902: begin
				q			<=			16'h000A;
		end
		32'h00009904: begin
				q			<=			16'hF097;
		end
		32'h00009906: begin
				q			<=			16'hFFFF;
		end
		32'h00009908: begin
				q			<=			16'h80E7;
		end
		32'h0000990A: begin
				q			<=			16'h2580;
		end
		32'h0000990C: begin
				q			<=			16'h0AE3;
		end
		32'h0000990E: begin
				q			<=			16'hBC05;
		end
		32'h00009910: begin
				q			<=			16'h5783;
		end
		32'h00009912: begin
				q			<=			16'h00C9;
		end
		32'h00009914: begin
				q			<=			16'hF793;
		end
		32'h00009916: begin
				q			<=			16'h0407;
		end
		32'h00009918: begin
				q			<=			16'h9663;
		end
		32'h0000991A: begin
				q			<=			16'hC807;
		end
		32'h0000991C: begin
				q			<=			16'h2083;
		end
		32'h0000991E: begin
				q			<=			16'h12C1;
		end
		32'h00009920: begin
				q			<=			16'h2403;
		end
		32'h00009922: begin
				q			<=			16'h1281;
		end
		32'h00009924: begin
				q			<=			16'h8513;
		end
		32'h00009926: begin
				q			<=			16'h000B;
		end
		32'h00009928: begin
				q			<=			16'h2483;
		end
		32'h0000992A: begin
				q			<=			16'h1241;
		end
		32'h0000992C: begin
				q			<=			16'h2903;
		end
		32'h0000992E: begin
				q			<=			16'h1201;
		end
		32'h00009930: begin
				q			<=			16'h2983;
		end
		32'h00009932: begin
				q			<=			16'h11C1;
		end
		32'h00009934: begin
				q			<=			16'h2A03;
		end
		32'h00009936: begin
				q			<=			16'h1181;
		end
		32'h00009938: begin
				q			<=			16'h2A83;
		end
		32'h0000993A: begin
				q			<=			16'h1141;
		end
		32'h0000993C: begin
				q			<=			16'h2B03;
		end
		32'h0000993E: begin
				q			<=			16'h1101;
		end
		32'h00009940: begin
				q			<=			16'h2B83;
		end
		32'h00009942: begin
				q			<=			16'h10C1;
		end
		32'h00009944: begin
				q			<=			16'h2C03;
		end
		32'h00009946: begin
				q			<=			16'h1081;
		end
		32'h00009948: begin
				q			<=			16'h2C83;
		end
		32'h0000994A: begin
				q			<=			16'h1041;
		end
		32'h0000994C: begin
				q			<=			16'h2D03;
		end
		32'h0000994E: begin
				q			<=			16'h1001;
		end
		32'h00009950: begin
				q			<=			16'h2D83;
		end
		32'h00009952: begin
				q			<=			16'h0FC1;
		end
		32'h00009954: begin
				q			<=			16'h0113;
		end
		32'h00009956: begin
				q			<=			16'h1301;
		end
		32'h00009958: begin
				q			<=			16'h8067;
		end
		32'h0000995A: begin
				q			<=			16'h0000;
		end
		32'h0000995C: begin
				q			<=			16'h8693;
		end
		32'h0000995E: begin
				q			<=			16'h0106;
		end
		32'h00009960: begin
				q			<=			16'h2223;
		end
		32'h00009962: begin
				q			<=			16'h0197;
		end
		32'h00009964: begin
				q			<=			16'h2423;
		end
		32'h00009966: begin
				q			<=			16'h04D1;
		end
		32'h00009968: begin
				q			<=			16'h2223;
		end
		32'h0000996A: begin
				q			<=			16'h04F1;
		end
		32'h0000996C: begin
				q			<=			16'h0713;
		end
		32'h0000996E: begin
				q			<=			16'h0087;
		end
		32'h00009970: begin
				q			<=			16'hD063;
		end
		32'h00009972: begin
				q			<=			16'h02FD;
		end
		32'h00009974: begin
				q			<=			16'h0613;
		end
		32'h00009976: begin
				q			<=			16'h0401;
		end
		32'h00009978: begin
				q			<=			16'h0593;
		end
		32'h0000997A: begin
				q			<=			16'h0009;
		end
		32'h0000997C: begin
				q			<=			16'h8513;
		end
		32'h0000997E: begin
				q			<=			16'h000A;
		end
		32'h00009980: begin
				q			<=			16'hF097;
		end
		32'h00009982: begin
				q			<=			16'hFFFF;
		end
		32'h00009984: begin
				q			<=			16'h80E7;
		end
		32'h00009986: begin
				q			<=			16'h1DC0;
		end
		32'h00009988: begin
				q			<=			16'h14E3;
		end
		32'h0000998A: begin
				q			<=			16'hF805;
		end
		32'h0000998C: begin
				q			<=			16'h0713;
		end
		32'h0000998E: begin
				q			<=			16'h000B;
		end
		32'h00009990: begin
				q			<=			16'h0413;
		end
		32'h00009992: begin
				q			<=			16'hFF04;
		end
		32'h00009994: begin
				q			<=			16'hF06F;
		end
		32'h00009996: begin
				q			<=			16'hF39F;
		end
		32'h00009998: begin
				q			<=			16'h2783;
		end
		32'h0000999A: begin
				q			<=			16'h0481;
		end
		32'h0000999C: begin
				q			<=			16'h8AE3;
		end
		32'h0000999E: begin
				q			<=			16'hF607;
		end
		32'h000099A0: begin
				q			<=			16'h0613;
		end
		32'h000099A2: begin
				q			<=			16'h0401;
		end
		32'h000099A4: begin
				q			<=			16'h0593;
		end
		32'h000099A6: begin
				q			<=			16'h0009;
		end
		32'h000099A8: begin
				q			<=			16'h8513;
		end
		32'h000099AA: begin
				q			<=			16'h000A;
		end
		32'h000099AC: begin
				q			<=			16'hF097;
		end
		32'h000099AE: begin
				q			<=			16'hFFFF;
		end
		32'h000099B0: begin
				q			<=			16'h80E7;
		end
		32'h000099B2: begin
				q			<=			16'h1B00;
		end
		32'h000099B4: begin
				q			<=			16'hF06F;
		end
		32'h000099B6: begin
				q			<=			16'hF5DF;
		end
		32'h000099B8: begin
				q			<=			16'h0000;
		end
		32'h000099BA: begin
				q			<=			16'h0000;
		end
		32'h000099BC: begin
				q			<=			16'h85B3;
		end
		32'h000099BE: begin
				q			<=			16'h02C5;
		end
		32'h000099C0: begin
				q			<=			16'h0113;
		end
		32'h000099C2: begin
				q			<=			16'hFF01;
		end
		32'h000099C4: begin
				q			<=			16'h2423;
		end
		32'h000099C6: begin
				q			<=			16'h0081;
		end
		32'h000099C8: begin
				q			<=			16'h2623;
		end
		32'h000099CA: begin
				q			<=			16'h0011;
		end
		32'h000099CC: begin
				q			<=			16'hD0EF;
		end
		32'h000099CE: begin
				q			<=			16'h9D5F;
		end
		32'h000099D0: begin
				q			<=			16'h0413;
		end
		32'h000099D2: begin
				q			<=			16'h0005;
		end
		32'h000099D4: begin
				q			<=			16'h0263;
		end
		32'h000099D6: begin
				q			<=			16'h0405;
		end
		32'h000099D8: begin
				q			<=			16'h2603;
		end
		32'h000099DA: begin
				q			<=			16'hFFC5;
		end
		32'h000099DC: begin
				q			<=			16'h0713;
		end
		32'h000099DE: begin
				q			<=			16'h0240;
		end
		32'h000099E0: begin
				q			<=			16'h7613;
		end
		32'h000099E2: begin
				q			<=			16'hFFC6;
		end
		32'h000099E4: begin
				q			<=			16'h0613;
		end
		32'h000099E6: begin
				q			<=			16'hFFC6;
		end
		32'h000099E8: begin
				q			<=			16'h6263;
		end
		32'h000099EA: begin
				q			<=			16'h06C7;
		end
		32'h000099EC: begin
				q			<=			16'h0693;
		end
		32'h000099EE: begin
				q			<=			16'h0130;
		end
		32'h000099F0: begin
				q			<=			16'h0793;
		end
		32'h000099F2: begin
				q			<=			16'h0005;
		end
		32'h000099F4: begin
				q			<=			16'hFC63;
		end
		32'h000099F6: begin
				q			<=			16'h00C6;
		end
		32'h000099F8: begin
				q			<=			16'h2023;
		end
		32'h000099FA: begin
				q			<=			16'h0005;
		end
		32'h000099FC: begin
				q			<=			16'h2223;
		end
		32'h000099FE: begin
				q			<=			16'h0005;
		end
		32'h00009A00: begin
				q			<=			16'h0793;
		end
		32'h00009A02: begin
				q			<=			16'h01B0;
		end
		32'h00009A04: begin
				q			<=			16'hE463;
		end
		32'h00009A06: begin
				q			<=			16'h02C7;
		end
		32'h00009A08: begin
				q			<=			16'h0793;
		end
		32'h00009A0A: begin
				q			<=			16'h0085;
		end
		32'h00009A0C: begin
				q			<=			16'hA023;
		end
		32'h00009A0E: begin
				q			<=			16'h0007;
		end
		32'h00009A10: begin
				q			<=			16'hA223;
		end
		32'h00009A12: begin
				q			<=			16'h0007;
		end
		32'h00009A14: begin
				q			<=			16'hA423;
		end
		32'h00009A16: begin
				q			<=			16'h0007;
		end
		32'h00009A18: begin
				q			<=			16'h0513;
		end
		32'h00009A1A: begin
				q			<=			16'h0004;
		end
		32'h00009A1C: begin
				q			<=			16'h2083;
		end
		32'h00009A1E: begin
				q			<=			16'h00C1;
		end
		32'h00009A20: begin
				q			<=			16'h2403;
		end
		32'h00009A22: begin
				q			<=			16'h0081;
		end
		32'h00009A24: begin
				q			<=			16'h0113;
		end
		32'h00009A26: begin
				q			<=			16'h0101;
		end
		32'h00009A28: begin
				q			<=			16'h8067;
		end
		32'h00009A2A: begin
				q			<=			16'h0000;
		end
		32'h00009A2C: begin
				q			<=			16'h2423;
		end
		32'h00009A2E: begin
				q			<=			16'h0005;
		end
		32'h00009A30: begin
				q			<=			16'h2623;
		end
		32'h00009A32: begin
				q			<=			16'h0005;
		end
		32'h00009A34: begin
				q			<=			16'h0793;
		end
		32'h00009A36: begin
				q			<=			16'h0105;
		end
		32'h00009A38: begin
				q			<=			16'h1AE3;
		end
		32'h00009A3A: begin
				q			<=			16'hFCE6;
		end
		32'h00009A3C: begin
				q			<=			16'h2823;
		end
		32'h00009A3E: begin
				q			<=			16'h0005;
		end
		32'h00009A40: begin
				q			<=			16'h0793;
		end
		32'h00009A42: begin
				q			<=			16'h0185;
		end
		32'h00009A44: begin
				q			<=			16'h2A23;
		end
		32'h00009A46: begin
				q			<=			16'h0005;
		end
		32'h00009A48: begin
				q			<=			16'hF06F;
		end
		32'h00009A4A: begin
				q			<=			16'hFC5F;
		end
		32'h00009A4C: begin
				q			<=			16'h0593;
		end
		32'h00009A4E: begin
				q			<=			16'h0000;
		end
		32'h00009A50: begin
				q			<=			16'h9097;
		end
		32'h00009A52: begin
				q			<=			16'hFFFF;
		end
		32'h00009A54: begin
				q			<=			16'h80E7;
		end
		32'h00009A56: begin
				q			<=			16'h1940;
		end
		32'h00009A58: begin
				q			<=			16'hF06F;
		end
		32'h00009A5A: begin
				q			<=			16'hFC1F;
		end
		32'h00009A5C: begin
				q			<=			16'h0000;
		end
		32'h00009A5E: begin
				q			<=			16'h0000;
		end
		32'h00009A60: begin
				q			<=			16'h0E63;
		end
		32'h00009A62: begin
				q			<=			16'h0606;
		end
		32'h00009A64: begin
				q			<=			16'h0113;
		end
		32'h00009A66: begin
				q			<=			16'hFF01;
		end
		32'h00009A68: begin
				q			<=			16'h6597;
		end
		32'h00009A6A: begin
				q			<=			16'h0000;
		end
		32'h00009A6C: begin
				q			<=			16'h8593;
		end
		32'h00009A6E: begin
				q			<=			16'h3745;
		end
		32'h00009A70: begin
				q			<=			16'h0513;
		end
		32'h00009A72: begin
				q			<=			16'h0006;
		end
		32'h00009A74: begin
				q			<=			16'h2423;
		end
		32'h00009A76: begin
				q			<=			16'h0081;
		end
		32'h00009A78: begin
				q			<=			16'h2623;
		end
		32'h00009A7A: begin
				q			<=			16'h0011;
		end
		32'h00009A7C: begin
				q			<=			16'h0413;
		end
		32'h00009A7E: begin
				q			<=			16'h0006;
		end
		32'h00009A80: begin
				q			<=			16'h1097;
		end
		32'h00009A82: begin
				q			<=			16'h0000;
		end
		32'h00009A84: begin
				q			<=			16'h80E7;
		end
		32'h00009A86: begin
				q			<=			16'h87C0;
		end
		32'h00009A88: begin
				q			<=			16'h0C63;
		end
		32'h00009A8A: begin
				q			<=			16'h0205;
		end
		32'h00009A8C: begin
				q			<=			16'h6597;
		end
		32'h00009A8E: begin
				q			<=			16'h0000;
		end
		32'h00009A90: begin
				q			<=			16'h8593;
		end
		32'h00009A92: begin
				q			<=			16'h34C5;
		end
		32'h00009A94: begin
				q			<=			16'h0513;
		end
		32'h00009A96: begin
				q			<=			16'h0004;
		end
		32'h00009A98: begin
				q			<=			16'h1097;
		end
		32'h00009A9A: begin
				q			<=			16'h0000;
		end
		32'h00009A9C: begin
				q			<=			16'h80E7;
		end
		32'h00009A9E: begin
				q			<=			16'h8640;
		end
		32'h00009AA0: begin
				q			<=			16'h0063;
		end
		32'h00009AA2: begin
				q			<=			16'h0205;
		end
		32'h00009AA4: begin
				q			<=			16'h6597;
		end
		32'h00009AA6: begin
				q			<=			16'h0000;
		end
		32'h00009AA8: begin
				q			<=			16'h8593;
		end
		32'h00009AAA: begin
				q			<=			16'h3045;
		end
		32'h00009AAC: begin
				q			<=			16'h0513;
		end
		32'h00009AAE: begin
				q			<=			16'h0004;
		end
		32'h00009AB0: begin
				q			<=			16'h1097;
		end
		32'h00009AB2: begin
				q			<=			16'h0000;
		end
		32'h00009AB4: begin
				q			<=			16'h80E7;
		end
		32'h00009AB6: begin
				q			<=			16'h84C0;
		end
		32'h00009AB8: begin
				q			<=			16'h0793;
		end
		32'h00009ABA: begin
				q			<=			16'h0000;
		end
		32'h00009ABC: begin
				q			<=			16'h1663;
		end
		32'h00009ABE: begin
				q			<=			16'h0005;
		end
		32'h00009AC0: begin
				q			<=			16'h6797;
		end
		32'h00009AC2: begin
				q			<=			16'h0000;
		end
		32'h00009AC4: begin
				q			<=			16'h8793;
		end
		32'h00009AC6: begin
				q			<=			16'h3187;
		end
		32'h00009AC8: begin
				q			<=			16'h2083;
		end
		32'h00009ACA: begin
				q			<=			16'h00C1;
		end
		32'h00009ACC: begin
				q			<=			16'h2403;
		end
		32'h00009ACE: begin
				q			<=			16'h0081;
		end
		32'h00009AD0: begin
				q			<=			16'h8513;
		end
		32'h00009AD2: begin
				q			<=			16'h0007;
		end
		32'h00009AD4: begin
				q			<=			16'h0113;
		end
		32'h00009AD6: begin
				q			<=			16'h0101;
		end
		32'h00009AD8: begin
				q			<=			16'h8067;
		end
		32'h00009ADA: begin
				q			<=			16'h0000;
		end
		32'h00009ADC: begin
				q			<=			16'h6797;
		end
		32'h00009ADE: begin
				q			<=			16'h0000;
		end
		32'h00009AE0: begin
				q			<=			16'h8793;
		end
		32'h00009AE2: begin
				q			<=			16'h2FC7;
		end
		32'h00009AE4: begin
				q			<=			16'h8513;
		end
		32'h00009AE6: begin
				q			<=			16'h0007;
		end
		32'h00009AE8: begin
				q			<=			16'h8067;
		end
		32'h00009AEA: begin
				q			<=			16'h0000;
		end
		32'h00009AEC: begin
				q			<=			16'h7797;
		end
		32'h00009AEE: begin
				q			<=			16'h0000;
		end
		32'h00009AF0: begin
				q			<=			16'h8793;
		end
		32'h00009AF2: begin
				q			<=			16'hDEC7;
		end
		32'h00009AF4: begin
				q			<=			16'hA783;
		end
		32'h00009AF6: begin
				q			<=			16'h0007;
		end
		32'h00009AF8: begin
				q			<=			16'hA783;
		end
		32'h00009AFA: begin
				q			<=			16'h0347;
		end
		32'h00009AFC: begin
				q			<=			16'h9663;
		end
		32'h00009AFE: begin
				q			<=			16'h0007;
		end
		32'h00009B00: begin
				q			<=			16'h7797;
		end
		32'h00009B02: begin
				q			<=			16'h0000;
		end
		32'h00009B04: begin
				q			<=			16'h8793;
		end
		32'h00009B06: begin
				q			<=			16'hC687;
		end
		32'h00009B08: begin
				q			<=			16'hC503;
		end
		32'h00009B0A: begin
				q			<=			16'h1287;
		end
		32'h00009B0C: begin
				q			<=			16'h8067;
		end
		32'h00009B0E: begin
				q			<=			16'h0000;
		end
		32'h00009B10: begin
				q			<=			16'h2503;
		end
		32'h00009B12: begin
				q			<=			16'h0EC5;
		end
		32'h00009B14: begin
				q			<=			16'h8067;
		end
		32'h00009B16: begin
				q			<=			16'h0000;
		end
		32'h00009B18: begin
				q			<=			16'h7797;
		end
		32'h00009B1A: begin
				q			<=			16'h0000;
		end
		32'h00009B1C: begin
				q			<=			16'h8793;
		end
		32'h00009B1E: begin
				q			<=			16'hDC07;
		end
		32'h00009B20: begin
				q			<=			16'hA783;
		end
		32'h00009B22: begin
				q			<=			16'h0007;
		end
		32'h00009B24: begin
				q			<=			16'hA783;
		end
		32'h00009B26: begin
				q			<=			16'h0347;
		end
		32'h00009B28: begin
				q			<=			16'h9663;
		end
		32'h00009B2A: begin
				q			<=			16'h0007;
		end
		32'h00009B2C: begin
				q			<=			16'h7797;
		end
		32'h00009B2E: begin
				q			<=			16'h0000;
		end
		32'h00009B30: begin
				q			<=			16'h8793;
		end
		32'h00009B32: begin
				q			<=			16'hC3C7;
		end
		32'h00009B34: begin
				q			<=			16'hA503;
		end
		32'h00009B36: begin
				q			<=			16'h0EC7;
		end
		32'h00009B38: begin
				q			<=			16'h8067;
		end
		32'h00009B3A: begin
				q			<=			16'h0000;
		end
		32'h00009B3C: begin
				q			<=			16'h7797;
		end
		32'h00009B3E: begin
				q			<=			16'h0000;
		end
		32'h00009B40: begin
				q			<=			16'h8793;
		end
		32'h00009B42: begin
				q			<=			16'hD9C7;
		end
		32'h00009B44: begin
				q			<=			16'h8613;
		end
		32'h00009B46: begin
				q			<=			16'h0005;
		end
		32'h00009B48: begin
				q			<=			16'h0593;
		end
		32'h00009B4A: begin
				q			<=			16'h0005;
		end
		32'h00009B4C: begin
				q			<=			16'hA503;
		end
		32'h00009B4E: begin
				q			<=			16'h0007;
		end
		32'h00009B50: begin
				q			<=			16'hF06F;
		end
		32'h00009B52: begin
				q			<=			16'hF11F;
		end
		32'h00009B54: begin
				q			<=			16'h0000;
		end
		32'h00009B56: begin
				q			<=			16'h0000;
		end
		32'h00009B58: begin
				q			<=			16'h7797;
		end
		32'h00009B5A: begin
				q			<=			16'h0000;
		end
		32'h00009B5C: begin
				q			<=			16'h8793;
		end
		32'h00009B5E: begin
				q			<=			16'hD807;
		end
		32'h00009B60: begin
				q			<=			16'hA783;
		end
		32'h00009B62: begin
				q			<=			16'h0007;
		end
		32'h00009B64: begin
				q			<=			16'hA783;
		end
		32'h00009B66: begin
				q			<=			16'h0347;
		end
		32'h00009B68: begin
				q			<=			16'h9663;
		end
		32'h00009B6A: begin
				q			<=			16'h0007;
		end
		32'h00009B6C: begin
				q			<=			16'h7797;
		end
		32'h00009B6E: begin
				q			<=			16'h0000;
		end
		32'h00009B70: begin
				q			<=			16'h8793;
		end
		32'h00009B72: begin
				q			<=			16'hBFC7;
		end
		32'h00009B74: begin
				q			<=			16'hA303;
		end
		32'h00009B76: begin
				q			<=			16'h0E47;
		end
		32'h00009B78: begin
				q			<=			16'h0067;
		end
		32'h00009B7A: begin
				q			<=			16'h0003;
		end
		32'h00009B7C: begin
				q			<=			16'h9A63;
		end
		32'h00009B7E: begin
				q			<=			16'h0205;
		end
		32'h00009B80: begin
				q			<=			16'h0113;
		end
		32'h00009B82: begin
				q			<=			16'hFF01;
		end
		32'h00009B84: begin
				q			<=			16'h0593;
		end
		32'h00009B86: begin
				q			<=			16'h00C1;
		end
		32'h00009B88: begin
				q			<=			16'h0513;
		end
		32'h00009B8A: begin
				q			<=			16'h0000;
		end
		32'h00009B8C: begin
				q			<=			16'h0E63;
		end
		32'h00009B8E: begin
				q			<=			16'h0006;
		end
		32'h00009B90: begin
				q			<=			16'h0513;
		end
		32'h00009B92: begin
				q			<=			16'hFFE0;
		end
		32'h00009B94: begin
				q			<=			16'h8A63;
		end
		32'h00009B96: begin
				q			<=			16'h0006;
		end
		32'h00009B98: begin
				q			<=			16'h4783;
		end
		32'h00009B9A: begin
				q			<=			16'h0006;
		end
		32'h00009B9C: begin
				q			<=			16'hA023;
		end
		32'h00009B9E: begin
				q			<=			16'h00F5;
		end
		32'h00009BA0: begin
				q			<=			16'h4503;
		end
		32'h00009BA2: begin
				q			<=			16'h0006;
		end
		32'h00009BA4: begin
				q			<=			16'h3533;
		end
		32'h00009BA6: begin
				q			<=			16'h00A0;
		end
		32'h00009BA8: begin
				q			<=			16'h0113;
		end
		32'h00009BAA: begin
				q			<=			16'h0101;
		end
		32'h00009BAC: begin
				q			<=			16'h8067;
		end
		32'h00009BAE: begin
				q			<=			16'h0000;
		end
		32'h00009BB0: begin
				q			<=			16'h0513;
		end
		32'h00009BB2: begin
				q			<=			16'h0000;
		end
		32'h00009BB4: begin
				q			<=			16'h0063;
		end
		32'h00009BB6: begin
				q			<=			16'h0206;
		end
		32'h00009BB8: begin
				q			<=			16'h0513;
		end
		32'h00009BBA: begin
				q			<=			16'hFFE0;
		end
		32'h00009BBC: begin
				q			<=			16'h8C63;
		end
		32'h00009BBE: begin
				q			<=			16'h0006;
		end
		32'h00009BC0: begin
				q			<=			16'h4783;
		end
		32'h00009BC2: begin
				q			<=			16'h0006;
		end
		32'h00009BC4: begin
				q			<=			16'hA023;
		end
		32'h00009BC6: begin
				q			<=			16'h00F5;
		end
		32'h00009BC8: begin
				q			<=			16'h4503;
		end
		32'h00009BCA: begin
				q			<=			16'h0006;
		end
		32'h00009BCC: begin
				q			<=			16'h3533;
		end
		32'h00009BCE: begin
				q			<=			16'h00A0;
		end
		32'h00009BD0: begin
				q			<=			16'h8067;
		end
		32'h00009BD2: begin
				q			<=			16'h0000;
		end
		32'h00009BD4: begin
				q			<=			16'h8067;
		end
		32'h00009BD6: begin
				q			<=			16'h0000;
		end
		32'h00009BD8: begin
				q			<=			16'h0000;
		end
		32'h00009BDA: begin
				q			<=			16'h0000;
		end
		32'h00009BDC: begin
				q			<=			16'h0733;
		end
		32'h00009BDE: begin
				q			<=			16'h00C5;
		end
		32'h00009BE0: begin
				q			<=			16'hE863;
		end
		32'h00009BE2: begin
				q			<=			16'h00A5;
		end
		32'h00009BE4: begin
				q			<=			16'h0793;
		end
		32'h00009BE6: begin
				q			<=			16'h0005;
		end
		32'h00009BE8: begin
				q			<=			16'h1A63;
		end
		32'h00009BEA: begin
				q			<=			16'h02F7;
		end
		32'h00009BEC: begin
				q			<=			16'h8067;
		end
		32'h00009BEE: begin
				q			<=			16'h0000;
		end
		32'h00009BF0: begin
				q			<=			16'h87B3;
		end
		32'h00009BF2: begin
				q			<=			16'h00C5;
		end
		32'h00009BF4: begin
				q			<=			16'h0633;
		end
		32'h00009BF6: begin
				q			<=			16'h40F6;
		end
		32'h00009BF8: begin
				q			<=			16'h76E3;
		end
		32'h00009BFA: begin
				q			<=			16'hFEF5;
		end
		32'h00009BFC: begin
				q			<=			16'h86B3;
		end
		32'h00009BFE: begin
				q			<=			16'h00C7;
		end
		32'h00009C00: begin
				q			<=			16'h9463;
		end
		32'h00009C02: begin
				q			<=			16'h0006;
		end
		32'h00009C04: begin
				q			<=			16'h8067;
		end
		32'h00009C06: begin
				q			<=			16'h0000;
		end
		32'h00009C08: begin
				q			<=			16'h8793;
		end
		32'h00009C0A: begin
				q			<=			16'hFFF7;
		end
		32'h00009C0C: begin
				q			<=			16'hC683;
		end
		32'h00009C0E: begin
				q			<=			16'h0007;
		end
		32'h00009C10: begin
				q			<=			16'h0713;
		end
		32'h00009C12: begin
				q			<=			16'hFFF7;
		end
		32'h00009C14: begin
				q			<=			16'h0023;
		end
		32'h00009C16: begin
				q			<=			16'h00D7;
		end
		32'h00009C18: begin
				q			<=			16'hF06F;
		end
		32'h00009C1A: begin
				q			<=			16'hFE5F;
		end
		32'h00009C1C: begin
				q			<=			16'h8593;
		end
		32'h00009C1E: begin
				q			<=			16'h0015;
		end
		32'h00009C20: begin
				q			<=			16'hC683;
		end
		32'h00009C22: begin
				q			<=			16'hFFF5;
		end
		32'h00009C24: begin
				q			<=			16'h8793;
		end
		32'h00009C26: begin
				q			<=			16'h0017;
		end
		32'h00009C28: begin
				q			<=			16'h8FA3;
		end
		32'h00009C2A: begin
				q			<=			16'hFED7;
		end
		32'h00009C2C: begin
				q			<=			16'hF06F;
		end
		32'h00009C2E: begin
				q			<=			16'hFBDF;
		end
		32'h00009C30: begin
				q			<=			16'h0000;
		end
		32'h00009C32: begin
				q			<=			16'h0000;
		end
		32'h00009C34: begin
				q			<=			16'h0113;
		end
		32'h00009C36: begin
				q			<=			16'hFC01;
		end
		32'h00009C38: begin
				q			<=			16'h2C23;
		end
		32'h00009C3A: begin
				q			<=			16'h0281;
		end
		32'h00009C3C: begin
				q			<=			16'h2E23;
		end
		32'h00009C3E: begin
				q			<=			16'h0211;
		end
		32'h00009C40: begin
				q			<=			16'h8413;
		end
		32'h00009C42: begin
				q			<=			16'h0005;
		end
		32'h00009C44: begin
				q			<=			16'h2A23;
		end
		32'h00009C46: begin
				q			<=			16'h0291;
		end
		32'h00009C48: begin
				q			<=			16'h2823;
		end
		32'h00009C4A: begin
				q			<=			16'h0321;
		end
		32'h00009C4C: begin
				q			<=			16'h2623;
		end
		32'h00009C4E: begin
				q			<=			16'h0331;
		end
		32'h00009C50: begin
				q			<=			16'h2423;
		end
		32'h00009C52: begin
				q			<=			16'h0341;
		end
		32'h00009C54: begin
				q			<=			16'h2223;
		end
		32'h00009C56: begin
				q			<=			16'h0351;
		end
		32'h00009C58: begin
				q			<=			16'h2023;
		end
		32'h00009C5A: begin
				q			<=			16'h0361;
		end
		32'h00009C5C: begin
				q			<=			16'h2E23;
		end
		32'h00009C5E: begin
				q			<=			16'h0171;
		end
		32'h00009C60: begin
				q			<=			16'h0593;
		end
		32'h00009C62: begin
				q			<=			16'h0006;
		end
		32'h00009C64: begin
				q			<=			16'h1863;
		end
		32'h00009C66: begin
				q			<=			16'h0204;
		end
		32'h00009C68: begin
				q			<=			16'h2403;
		end
		32'h00009C6A: begin
				q			<=			16'h0381;
		end
		32'h00009C6C: begin
				q			<=			16'h2083;
		end
		32'h00009C6E: begin
				q			<=			16'h03C1;
		end
		32'h00009C70: begin
				q			<=			16'h2483;
		end
		32'h00009C72: begin
				q			<=			16'h0341;
		end
		32'h00009C74: begin
				q			<=			16'h2903;
		end
		32'h00009C76: begin
				q			<=			16'h0301;
		end
		32'h00009C78: begin
				q			<=			16'h2983;
		end
		32'h00009C7A: begin
				q			<=			16'h02C1;
		end
		32'h00009C7C: begin
				q			<=			16'h2A03;
		end
		32'h00009C7E: begin
				q			<=			16'h0281;
		end
		32'h00009C80: begin
				q			<=			16'h2A83;
		end
		32'h00009C82: begin
				q			<=			16'h0241;
		end
		32'h00009C84: begin
				q			<=			16'h2B03;
		end
		32'h00009C86: begin
				q			<=			16'h0201;
		end
		32'h00009C88: begin
				q			<=			16'h2B83;
		end
		32'h00009C8A: begin
				q			<=			16'h01C1;
		end
		32'h00009C8C: begin
				q			<=			16'h0113;
		end
		32'h00009C8E: begin
				q			<=			16'h0401;
		end
		32'h00009C90: begin
				q			<=			16'hD06F;
		end
		32'h00009C92: begin
				q			<=			16'hF10F;
		end
		32'h00009C94: begin
				q			<=			16'h0A93;
		end
		32'h00009C96: begin
				q			<=			16'h0005;
		end
		32'h00009C98: begin
				q			<=			16'h2623;
		end
		32'h00009C9A: begin
				q			<=			16'h00C1;
		end
		32'h00009C9C: begin
				q			<=			16'hD0EF;
		end
		32'h00009C9E: begin
				q			<=			16'hDE5F;
		end
		32'h00009CA0: begin
				q			<=			16'h2583;
		end
		32'h00009CA2: begin
				q			<=			16'h00C1;
		end
		32'h00009CA4: begin
				q			<=			16'h2683;
		end
		32'h00009CA6: begin
				q			<=			16'hFFC4;
		end
		32'h00009CA8: begin
				q			<=			16'h0793;
		end
		32'h00009CAA: begin
				q			<=			16'h0160;
		end
		32'h00009CAC: begin
				q			<=			16'h8993;
		end
		32'h00009CAE: begin
				q			<=			16'h00B5;
		end
		32'h00009CB0: begin
				q			<=			16'h0B93;
		end
		32'h00009CB2: begin
				q			<=			16'hFF84;
		end
		32'h00009CB4: begin
				q			<=			16'hF913;
		end
		32'h00009CB6: begin
				q			<=			16'hFFC6;
		end
		32'h00009CB8: begin
				q			<=			16'hF463;
		end
		32'h00009CBA: begin
				q			<=			16'h0537;
		end
		32'h00009CBC: begin
				q			<=			16'hFB13;
		end
		32'h00009CBE: begin
				q			<=			16'hFF89;
		end
		32'h00009CC0: begin
				q			<=			16'h5263;
		end
		32'h00009CC2: begin
				q			<=			16'h040B;
		end
		32'h00009CC4: begin
				q			<=			16'h0793;
		end
		32'h00009CC6: begin
				q			<=			16'h00C0;
		end
		32'h00009CC8: begin
				q			<=			16'hA023;
		end
		32'h00009CCA: begin
				q			<=			16'h00FA;
		end
		32'h00009CCC: begin
				q			<=			16'h0A13;
		end
		32'h00009CCE: begin
				q			<=			16'h0000;
		end
		32'h00009CD0: begin
				q			<=			16'h2083;
		end
		32'h00009CD2: begin
				q			<=			16'h03C1;
		end
		32'h00009CD4: begin
				q			<=			16'h2403;
		end
		32'h00009CD6: begin
				q			<=			16'h0381;
		end
		32'h00009CD8: begin
				q			<=			16'h0513;
		end
		32'h00009CDA: begin
				q			<=			16'h000A;
		end
		32'h00009CDC: begin
				q			<=			16'h2483;
		end
		32'h00009CDE: begin
				q			<=			16'h0341;
		end
		32'h00009CE0: begin
				q			<=			16'h2903;
		end
		32'h00009CE2: begin
				q			<=			16'h0301;
		end
		32'h00009CE4: begin
				q			<=			16'h2983;
		end
		32'h00009CE6: begin
				q			<=			16'h02C1;
		end
		32'h00009CE8: begin
				q			<=			16'h2A03;
		end
		32'h00009CEA: begin
				q			<=			16'h0281;
		end
		32'h00009CEC: begin
				q			<=			16'h2A83;
		end
		32'h00009CEE: begin
				q			<=			16'h0241;
		end
		32'h00009CF0: begin
				q			<=			16'h2B03;
		end
		32'h00009CF2: begin
				q			<=			16'h0201;
		end
		32'h00009CF4: begin
				q			<=			16'h2B83;
		end
		32'h00009CF6: begin
				q			<=			16'h01C1;
		end
		32'h00009CF8: begin
				q			<=			16'h0113;
		end
		32'h00009CFA: begin
				q			<=			16'h0401;
		end
		32'h00009CFC: begin
				q			<=			16'h8067;
		end
		32'h00009CFE: begin
				q			<=			16'h0000;
		end
		32'h00009D00: begin
				q			<=			16'h0B13;
		end
		32'h00009D02: begin
				q			<=			16'h0100;
		end
		32'h00009D04: begin
				q			<=			16'h60E3;
		end
		32'h00009D06: begin
				q			<=			16'hFCBB;
		end
		32'h00009D08: begin
				q			<=			16'h5863;
		end
		32'h00009D0A: begin
				q			<=			16'h4769;
		end
		32'h00009D0C: begin
				q			<=			16'h6717;
		end
		32'h00009D0E: begin
				q			<=			16'h0000;
		end
		32'h00009D10: begin
				q			<=			16'h0713;
		end
		32'h00009D12: begin
				q			<=			16'h6547;
		end
		32'h00009D14: begin
				q			<=			16'h2603;
		end
		32'h00009D16: begin
				q			<=			16'h0087;
		end
		32'h00009D18: begin
				q			<=			16'h87B3;
		end
		32'h00009D1A: begin
				q			<=			16'h012B;
		end
		32'h00009D1C: begin
				q			<=			16'hA703;
		end
		32'h00009D1E: begin
				q			<=			16'h0047;
		end
		32'h00009D20: begin
				q			<=			16'h0C63;
		end
		32'h00009D22: begin
				q			<=			16'h00F6;
		end
		32'h00009D24: begin
				q			<=			16'h7513;
		end
		32'h00009D26: begin
				q			<=			16'hFFE7;
		end
		32'h00009D28: begin
				q			<=			16'h8533;
		end
		32'h00009D2A: begin
				q			<=			16'h00A7;
		end
		32'h00009D2C: begin
				q			<=			16'h2503;
		end
		32'h00009D2E: begin
				q			<=			16'h0045;
		end
		32'h00009D30: begin
				q			<=			16'h7513;
		end
		32'h00009D32: begin
				q			<=			16'h0015;
		end
		32'h00009D34: begin
				q			<=			16'h1263;
		end
		32'h00009D36: begin
				q			<=			16'h0C05;
		end
		32'h00009D38: begin
				q			<=			16'h7713;
		end
		32'h00009D3A: begin
				q			<=			16'hFFC7;
		end
		32'h00009D3C: begin
				q			<=			16'h09B3;
		end
		32'h00009D3E: begin
				q			<=			16'h00E9;
		end
		32'h00009D40: begin
				q			<=			16'h1463;
		end
		32'h00009D42: begin
				q			<=			16'h04F6;
		end
		32'h00009D44: begin
				q			<=			16'h0513;
		end
		32'h00009D46: begin
				q			<=			16'h010B;
		end
		32'h00009D48: begin
				q			<=			16'hCC63;
		end
		32'h00009D4A: begin
				q			<=			16'h0AA9;
		end
		32'h00009D4C: begin
				q			<=			16'h8BB3;
		end
		32'h00009D4E: begin
				q			<=			16'h016B;
		end
		32'h00009D50: begin
				q			<=			16'h89B3;
		end
		32'h00009D52: begin
				q			<=			16'h4169;
		end
		32'h00009D54: begin
				q			<=			16'h6797;
		end
		32'h00009D56: begin
				q			<=			16'h0000;
		end
		32'h00009D58: begin
				q			<=			16'hAA23;
		end
		32'h00009D5A: begin
				q			<=			16'h6177;
		end
		32'h00009D5C: begin
				q			<=			16'hE993;
		end
		32'h00009D5E: begin
				q			<=			16'h0019;
		end
		32'h00009D60: begin
				q			<=			16'hA223;
		end
		32'h00009D62: begin
				q			<=			16'h013B;
		end
		32'h00009D64: begin
				q			<=			16'h2983;
		end
		32'h00009D66: begin
				q			<=			16'hFFC4;
		end
		32'h00009D68: begin
				q			<=			16'h8513;
		end
		32'h00009D6A: begin
				q			<=			16'h000A;
		end
		32'h00009D6C: begin
				q			<=			16'h0A13;
		end
		32'h00009D6E: begin
				q			<=			16'h0004;
		end
		32'h00009D70: begin
				q			<=			16'hF993;
		end
		32'h00009D72: begin
				q			<=			16'h0019;
		end
		32'h00009D74: begin
				q			<=			16'hE9B3;
		end
		32'h00009D76: begin
				q			<=			16'h0169;
		end
		32'h00009D78: begin
				q			<=			16'h2E23;
		end
		32'h00009D7A: begin
				q			<=			16'hFF34;
		end
		32'h00009D7C: begin
				q			<=			16'hE097;
		end
		32'h00009D7E: begin
				q			<=			16'hFFFF;
		end
		32'h00009D80: begin
				q			<=			16'h80E7;
		end
		32'h00009D82: begin
				q			<=			16'hD080;
		end
		32'h00009D84: begin
				q			<=			16'hF06F;
		end
		32'h00009D86: begin
				q			<=			16'hF4DF;
		end
		32'h00009D88: begin
				q			<=			16'hCC63;
		end
		32'h00009D8A: begin
				q			<=			16'h0769;
		end
		32'h00009D8C: begin
				q			<=			16'hA703;
		end
		32'h00009D8E: begin
				q			<=			16'h00C7;
		end
		32'h00009D90: begin
				q			<=			16'hA783;
		end
		32'h00009D92: begin
				q			<=			16'h0087;
		end
		32'h00009D94: begin
				q			<=			16'hA623;
		end
		32'h00009D96: begin
				q			<=			16'h00E7;
		end
		32'h00009D98: begin
				q			<=			16'h2423;
		end
		32'h00009D9A: begin
				q			<=			16'h00F7;
		end
		32'h00009D9C: begin
				q			<=			16'hA703;
		end
		32'h00009D9E: begin
				q			<=			16'h004B;
		end
		32'h00009DA0: begin
				q			<=			16'h86B3;
		end
		32'h00009DA2: begin
				q			<=			16'h4169;
		end
		32'h00009DA4: begin
				q			<=			16'h0613;
		end
		32'h00009DA6: begin
				q			<=			16'h00F0;
		end
		32'h00009DA8: begin
				q			<=			16'h7713;
		end
		32'h00009DAA: begin
				q			<=			16'h0017;
		end
		32'h00009DAC: begin
				q			<=			16'h87B3;
		end
		32'h00009DAE: begin
				q			<=			16'h013B;
		end
		32'h00009DB0: begin
				q			<=			16'h7863;
		end
		32'h00009DB2: begin
				q			<=			16'h3CD6;
		end
		32'h00009DB4: begin
				q			<=			16'h69B3;
		end
		32'h00009DB6: begin
				q			<=			16'h00EB;
		end
		32'h00009DB8: begin
				q			<=			16'hA223;
		end
		32'h00009DBA: begin
				q			<=			16'h013B;
		end
		32'h00009DBC: begin
				q			<=			16'h85B3;
		end
		32'h00009DBE: begin
				q			<=			16'h016B;
		end
		32'h00009DC0: begin
				q			<=			16'hE693;
		end
		32'h00009DC2: begin
				q			<=			16'h0016;
		end
		32'h00009DC4: begin
				q			<=			16'hA223;
		end
		32'h00009DC6: begin
				q			<=			16'h00D5;
		end
		32'h00009DC8: begin
				q			<=			16'hA703;
		end
		32'h00009DCA: begin
				q			<=			16'h0047;
		end
		32'h00009DCC: begin
				q			<=			16'h8593;
		end
		32'h00009DCE: begin
				q			<=			16'h0085;
		end
		32'h00009DD0: begin
				q			<=			16'h8513;
		end
		32'h00009DD2: begin
				q			<=			16'h000A;
		end
		32'h00009DD4: begin
				q			<=			16'h6713;
		end
		32'h00009DD6: begin
				q			<=			16'h0017;
		end
		32'h00009DD8: begin
				q			<=			16'hA223;
		end
		32'h00009DDA: begin
				q			<=			16'h00E7;
		end
		32'h00009DDC: begin
				q			<=			16'hB097;
		end
		32'h00009DDE: begin
				q			<=			16'hFFFF;
		end
		32'h00009DE0: begin
				q			<=			16'h80E7;
		end
		32'h00009DE2: begin
				q			<=			16'h1940;
		end
		32'h00009DE4: begin
				q			<=			16'h8513;
		end
		32'h00009DE6: begin
				q			<=			16'h000A;
		end
		32'h00009DE8: begin
				q			<=			16'hE097;
		end
		32'h00009DEA: begin
				q			<=			16'hFFFF;
		end
		32'h00009DEC: begin
				q			<=			16'h80E7;
		end
		32'h00009DEE: begin
				q			<=			16'hC9C0;
		end
		32'h00009DF0: begin
				q			<=			16'h8A13;
		end
		32'h00009DF2: begin
				q			<=			16'h008B;
		end
		32'h00009DF4: begin
				q			<=			16'hF06F;
		end
		32'h00009DF6: begin
				q			<=			16'hEDDF;
		end
		32'h00009DF8: begin
				q			<=			16'h0713;
		end
		32'h00009DFA: begin
				q			<=			16'h0000;
		end
		32'h00009DFC: begin
				q			<=			16'h0793;
		end
		32'h00009DFE: begin
				q			<=			16'h0000;
		end
		32'h00009E00: begin
				q			<=			16'hF693;
		end
		32'h00009E02: begin
				q			<=			16'h0016;
		end
		32'h00009E04: begin
				q			<=			16'h9663;
		end
		32'h00009E06: begin
				q			<=			16'h2806;
		end
		32'h00009E08: begin
				q			<=			16'h2483;
		end
		32'h00009E0A: begin
				q			<=			16'hFF84;
		end
		32'h00009E0C: begin
				q			<=			16'h84B3;
		end
		32'h00009E0E: begin
				q			<=			16'h409B;
		end
		32'h00009E10: begin
				q			<=			16'hAA03;
		end
		32'h00009E12: begin
				q			<=			16'h0044;
		end
		32'h00009E14: begin
				q			<=			16'h7A13;
		end
		32'h00009E16: begin
				q			<=			16'hFFCA;
		end
		32'h00009E18: begin
				q			<=			16'h0A33;
		end
		32'h00009E1A: begin
				q			<=			16'h012A;
		end
		32'h00009E1C: begin
				q			<=			16'h8063;
		end
		32'h00009E1E: begin
				q			<=			16'h1C07;
		end
		32'h00009E20: begin
				q			<=			16'h09B3;
		end
		32'h00009E22: begin
				q			<=			16'h0147;
		end
		32'h00009E24: begin
				q			<=			16'h1A63;
		end
		32'h00009E26: begin
				q			<=			16'h0EF6;
		end
		32'h00009E28: begin
				q			<=			16'h0793;
		end
		32'h00009E2A: begin
				q			<=			16'h010B;
		end
		32'h00009E2C: begin
				q			<=			16'hC863;
		end
		32'h00009E2E: begin
				q			<=			16'h1AF9;
		end
		32'h00009E30: begin
				q			<=			16'hA703;
		end
		32'h00009E32: begin
				q			<=			16'h0084;
		end
		32'h00009E34: begin
				q			<=			16'hA783;
		end
		32'h00009E36: begin
				q			<=			16'h00C4;
		end
		32'h00009E38: begin
				q			<=			16'h0613;
		end
		32'h00009E3A: begin
				q			<=			16'hFFC9;
		end
		32'h00009E3C: begin
				q			<=			16'h8A13;
		end
		32'h00009E3E: begin
				q			<=			16'h0084;
		end
		32'h00009E40: begin
				q			<=			16'h2623;
		end
		32'h00009E42: begin
				q			<=			16'h00F7;
		end
		32'h00009E44: begin
				q			<=			16'hA423;
		end
		32'h00009E46: begin
				q			<=			16'h00E7;
		end
		32'h00009E48: begin
				q			<=			16'h0713;
		end
		32'h00009E4A: begin
				q			<=			16'h0240;
		end
		32'h00009E4C: begin
				q			<=			16'h6E63;
		end
		32'h00009E4E: begin
				q			<=			16'h0AC7;
		end
		32'h00009E50: begin
				q			<=			16'h0693;
		end
		32'h00009E52: begin
				q			<=			16'h0130;
		end
		32'h00009E54: begin
				q			<=			16'h0793;
		end
		32'h00009E56: begin
				q			<=			16'h000A;
		end
		32'h00009E58: begin
				q			<=			16'hF263;
		end
		32'h00009E5A: begin
				q			<=			16'h02C6;
		end
		32'h00009E5C: begin
				q			<=			16'h2783;
		end
		32'h00009E5E: begin
				q			<=			16'h0004;
		end
		32'h00009E60: begin
				q			<=			16'hA423;
		end
		32'h00009E62: begin
				q			<=			16'h00F4;
		end
		32'h00009E64: begin
				q			<=			16'h2783;
		end
		32'h00009E66: begin
				q			<=			16'h0044;
		end
		32'h00009E68: begin
				q			<=			16'hA623;
		end
		32'h00009E6A: begin
				q			<=			16'h00F4;
		end
		32'h00009E6C: begin
				q			<=			16'h0793;
		end
		32'h00009E6E: begin
				q			<=			16'h01B0;
		end
		32'h00009E70: begin
				q			<=			16'hEE63;
		end
		32'h00009E72: begin
				q			<=			16'h04C7;
		end
		32'h00009E74: begin
				q			<=			16'h0413;
		end
		32'h00009E76: begin
				q			<=			16'h0084;
		end
		32'h00009E78: begin
				q			<=			16'h8793;
		end
		32'h00009E7A: begin
				q			<=			16'h0104;
		end
		32'h00009E7C: begin
				q			<=			16'h2703;
		end
		32'h00009E7E: begin
				q			<=			16'h0004;
		end
		32'h00009E80: begin
				q			<=			16'hA023;
		end
		32'h00009E82: begin
				q			<=			16'h00E7;
		end
		32'h00009E84: begin
				q			<=			16'h2703;
		end
		32'h00009E86: begin
				q			<=			16'h0044;
		end
		32'h00009E88: begin
				q			<=			16'hA223;
		end
		32'h00009E8A: begin
				q			<=			16'h00E7;
		end
		32'h00009E8C: begin
				q			<=			16'h2703;
		end
		32'h00009E8E: begin
				q			<=			16'h0084;
		end
		32'h00009E90: begin
				q			<=			16'hA423;
		end
		32'h00009E92: begin
				q			<=			16'h00E7;
		end
		32'h00009E94: begin
				q			<=			16'h87B3;
		end
		32'h00009E96: begin
				q			<=			16'h0164;
		end
		32'h00009E98: begin
				q			<=			16'h89B3;
		end
		32'h00009E9A: begin
				q			<=			16'h4169;
		end
		32'h00009E9C: begin
				q			<=			16'h6717;
		end
		32'h00009E9E: begin
				q			<=			16'h0000;
		end
		32'h00009EA0: begin
				q			<=			16'h2623;
		end
		32'h00009EA2: begin
				q			<=			16'h4CF7;
		end
		32'h00009EA4: begin
				q			<=			16'hE993;
		end
		32'h00009EA6: begin
				q			<=			16'h0019;
		end
		32'h00009EA8: begin
				q			<=			16'hA223;
		end
		32'h00009EAA: begin
				q			<=			16'h0137;
		end
		32'h00009EAC: begin
				q			<=			16'hA783;
		end
		32'h00009EAE: begin
				q			<=			16'h0044;
		end
		32'h00009EB0: begin
				q			<=			16'hF793;
		end
		32'h00009EB2: begin
				q			<=			16'h0017;
		end
		32'h00009EB4: begin
				q			<=			16'hE9B3;
		end
		32'h00009EB6: begin
				q			<=			16'h0167;
		end
		32'h00009EB8: begin
				q			<=			16'hA223;
		end
		32'h00009EBA: begin
				q			<=			16'h0134;
		end
		32'h00009EBC: begin
				q			<=			16'h8513;
		end
		32'h00009EBE: begin
				q			<=			16'h000A;
		end
		32'h00009EC0: begin
				q			<=			16'hE097;
		end
		32'h00009EC2: begin
				q			<=			16'hFFFF;
		end
		32'h00009EC4: begin
				q			<=			16'h80E7;
		end
		32'h00009EC6: begin
				q			<=			16'hBC40;
		end
		32'h00009EC8: begin
				q			<=			16'hF06F;
		end
		32'h00009ECA: begin
				q			<=			16'hE09F;
		end
		32'h00009ECC: begin
				q			<=			16'h2783;
		end
		32'h00009ECE: begin
				q			<=			16'h0084;
		end
		32'h00009ED0: begin
				q			<=			16'hA823;
		end
		32'h00009ED2: begin
				q			<=			16'h00F4;
		end
		32'h00009ED4: begin
				q			<=			16'h2783;
		end
		32'h00009ED6: begin
				q			<=			16'h00C4;
		end
		32'h00009ED8: begin
				q			<=			16'hAA23;
		end
		32'h00009EDA: begin
				q			<=			16'h00F4;
		end
		32'h00009EDC: begin
				q			<=			16'h0863;
		end
		32'h00009EDE: begin
				q			<=			16'h00E6;
		end
		32'h00009EE0: begin
				q			<=			16'h0413;
		end
		32'h00009EE2: begin
				q			<=			16'h0104;
		end
		32'h00009EE4: begin
				q			<=			16'h8793;
		end
		32'h00009EE6: begin
				q			<=			16'h0184;
		end
		32'h00009EE8: begin
				q			<=			16'hF06F;
		end
		32'h00009EEA: begin
				q			<=			16'hF95F;
		end
		32'h00009EEC: begin
				q			<=			16'h2783;
		end
		32'h00009EEE: begin
				q			<=			16'h0104;
		end
		32'h00009EF0: begin
				q			<=			16'h0413;
		end
		32'h00009EF2: begin
				q			<=			16'h0184;
		end
		32'h00009EF4: begin
				q			<=			16'hAC23;
		end
		32'h00009EF6: begin
				q			<=			16'h00F4;
		end
		32'h00009EF8: begin
				q			<=			16'h2703;
		end
		32'h00009EFA: begin
				q			<=			16'hFFC4;
		end
		32'h00009EFC: begin
				q			<=			16'h8793;
		end
		32'h00009EFE: begin
				q			<=			16'h0204;
		end
		32'h00009F00: begin
				q			<=			16'hAE23;
		end
		32'h00009F02: begin
				q			<=			16'h00E4;
		end
		32'h00009F04: begin
				q			<=			16'hF06F;
		end
		32'h00009F06: begin
				q			<=			16'hF79F;
		end
		32'h00009F08: begin
				q			<=			16'h0593;
		end
		32'h00009F0A: begin
				q			<=			16'h0004;
		end
		32'h00009F0C: begin
				q			<=			16'h0513;
		end
		32'h00009F0E: begin
				q			<=			16'h000A;
		end
		32'h00009F10: begin
				q			<=			16'hF0EF;
		end
		32'h00009F12: begin
				q			<=			16'hCCDF;
		end
		32'h00009F14: begin
				q			<=			16'hF06F;
		end
		32'h00009F16: begin
				q			<=			16'hF81F;
		end
		32'h00009F18: begin
				q			<=			16'hC263;
		end
		32'h00009F1A: begin
				q			<=			16'h0D69;
		end
		32'h00009F1C: begin
				q			<=			16'hA703;
		end
		32'h00009F1E: begin
				q			<=			16'h00C7;
		end
		32'h00009F20: begin
				q			<=			16'hA783;
		end
		32'h00009F22: begin
				q			<=			16'h0087;
		end
		32'h00009F24: begin
				q			<=			16'h0613;
		end
		32'h00009F26: begin
				q			<=			16'hFFC9;
		end
		32'h00009F28: begin
				q			<=			16'h8513;
		end
		32'h00009F2A: begin
				q			<=			16'h0084;
		end
		32'h00009F2C: begin
				q			<=			16'hA623;
		end
		32'h00009F2E: begin
				q			<=			16'h00E7;
		end
		32'h00009F30: begin
				q			<=			16'h2423;
		end
		32'h00009F32: begin
				q			<=			16'h00F7;
		end
		32'h00009F34: begin
				q			<=			16'hA703;
		end
		32'h00009F36: begin
				q			<=			16'h0084;
		end
		32'h00009F38: begin
				q			<=			16'hA783;
		end
		32'h00009F3A: begin
				q			<=			16'h00C4;
		end
		32'h00009F3C: begin
				q			<=			16'h2623;
		end
		32'h00009F3E: begin
				q			<=			16'h00F7;
		end
		32'h00009F40: begin
				q			<=			16'hA423;
		end
		32'h00009F42: begin
				q			<=			16'h00E7;
		end
		32'h00009F44: begin
				q			<=			16'h0793;
		end
		32'h00009F46: begin
				q			<=			16'h0240;
		end
		32'h00009F48: begin
				q			<=			16'hE463;
		end
		32'h00009F4A: begin
				q			<=			16'h08C7;
		end
		32'h00009F4C: begin
				q			<=			16'h0713;
		end
		32'h00009F4E: begin
				q			<=			16'h0130;
		end
		32'h00009F50: begin
				q			<=			16'h7263;
		end
		32'h00009F52: begin
				q			<=			16'h02C7;
		end
		32'h00009F54: begin
				q			<=			16'h2703;
		end
		32'h00009F56: begin
				q			<=			16'h0004;
		end
		32'h00009F58: begin
				q			<=			16'hA423;
		end
		32'h00009F5A: begin
				q			<=			16'h00E4;
		end
		32'h00009F5C: begin
				q			<=			16'h2703;
		end
		32'h00009F5E: begin
				q			<=			16'h0044;
		end
		32'h00009F60: begin
				q			<=			16'hA623;
		end
		32'h00009F62: begin
				q			<=			16'h00E4;
		end
		32'h00009F64: begin
				q			<=			16'h0713;
		end
		32'h00009F66: begin
				q			<=			16'h01B0;
		end
		32'h00009F68: begin
				q			<=			16'h6663;
		end
		32'h00009F6A: begin
				q			<=			16'h02C7;
		end
		32'h00009F6C: begin
				q			<=			16'h0413;
		end
		32'h00009F6E: begin
				q			<=			16'h0084;
		end
		32'h00009F70: begin
				q			<=			16'h8513;
		end
		32'h00009F72: begin
				q			<=			16'h0104;
		end
		32'h00009F74: begin
				q			<=			16'h2783;
		end
		32'h00009F76: begin
				q			<=			16'h0004;
		end
		32'h00009F78: begin
				q			<=			16'h2023;
		end
		32'h00009F7A: begin
				q			<=			16'h00F5;
		end
		32'h00009F7C: begin
				q			<=			16'h2783;
		end
		32'h00009F7E: begin
				q			<=			16'h0044;
		end
		32'h00009F80: begin
				q			<=			16'h2223;
		end
		32'h00009F82: begin
				q			<=			16'h00F5;
		end
		32'h00009F84: begin
				q			<=			16'h2783;
		end
		32'h00009F86: begin
				q			<=			16'h0084;
		end
		32'h00009F88: begin
				q			<=			16'h2423;
		end
		32'h00009F8A: begin
				q			<=			16'h00F5;
		end
		32'h00009F8C: begin
				q			<=			16'h8B93;
		end
		32'h00009F8E: begin
				q			<=			16'h0004;
		end
		32'h00009F90: begin
				q			<=			16'hF06F;
		end
		32'h00009F92: begin
				q			<=			16'hE0DF;
		end
		32'h00009F94: begin
				q			<=			16'h2703;
		end
		32'h00009F96: begin
				q			<=			16'h0084;
		end
		32'h00009F98: begin
				q			<=			16'hA823;
		end
		32'h00009F9A: begin
				q			<=			16'h00E4;
		end
		32'h00009F9C: begin
				q			<=			16'h2703;
		end
		32'h00009F9E: begin
				q			<=			16'h00C4;
		end
		32'h00009FA0: begin
				q			<=			16'hAA23;
		end
		32'h00009FA2: begin
				q			<=			16'h00E4;
		end
		32'h00009FA4: begin
				q			<=			16'h0863;
		end
		32'h00009FA6: begin
				q			<=			16'h00F6;
		end
		32'h00009FA8: begin
				q			<=			16'h0413;
		end
		32'h00009FAA: begin
				q			<=			16'h0104;
		end
		32'h00009FAC: begin
				q			<=			16'h8513;
		end
		32'h00009FAE: begin
				q			<=			16'h0184;
		end
		32'h00009FB0: begin
				q			<=			16'hF06F;
		end
		32'h00009FB2: begin
				q			<=			16'hFC5F;
		end
		32'h00009FB4: begin
				q			<=			16'h2783;
		end
		32'h00009FB6: begin
				q			<=			16'h0104;
		end
		32'h00009FB8: begin
				q			<=			16'h8513;
		end
		32'h00009FBA: begin
				q			<=			16'h0204;
		end
		32'h00009FBC: begin
				q			<=			16'h0413;
		end
		32'h00009FBE: begin
				q			<=			16'h0184;
		end
		32'h00009FC0: begin
				q			<=			16'hAC23;
		end
		32'h00009FC2: begin
				q			<=			16'h00F4;
		end
		32'h00009FC4: begin
				q			<=			16'h2783;
		end
		32'h00009FC6: begin
				q			<=			16'hFFC4;
		end
		32'h00009FC8: begin
				q			<=			16'hAE23;
		end
		32'h00009FCA: begin
				q			<=			16'h00F4;
		end
		32'h00009FCC: begin
				q			<=			16'hF06F;
		end
		32'h00009FCE: begin
				q			<=			16'hFA9F;
		end
		32'h00009FD0: begin
				q			<=			16'h0593;
		end
		32'h00009FD2: begin
				q			<=			16'h0004;
		end
		32'h00009FD4: begin
				q			<=			16'hF0EF;
		end
		32'h00009FD6: begin
				q			<=			16'hC09F;
		end
		32'h00009FD8: begin
				q			<=			16'hF06F;
		end
		32'h00009FDA: begin
				q			<=			16'hFB5F;
		end
		32'h00009FDC: begin
				q			<=			16'h4A63;
		end
		32'h00009FDE: begin
				q			<=			16'h0B6A;
		end
		32'h00009FE0: begin
				q			<=			16'hA783;
		end
		32'h00009FE2: begin
				q			<=			16'h00C4;
		end
		32'h00009FE4: begin
				q			<=			16'hA703;
		end
		32'h00009FE6: begin
				q			<=			16'h0084;
		end
		32'h00009FE8: begin
				q			<=			16'h0613;
		end
		32'h00009FEA: begin
				q			<=			16'hFFC9;
		end
		32'h00009FEC: begin
				q			<=			16'h8513;
		end
		32'h00009FEE: begin
				q			<=			16'h0084;
		end
		32'h00009FF0: begin
				q			<=			16'h2623;
		end
		32'h00009FF2: begin
				q			<=			16'h00F7;
		end
		32'h00009FF4: begin
				q			<=			16'hA423;
		end
		32'h00009FF6: begin
				q			<=			16'h00E7;
		end
		32'h00009FF8: begin
				q			<=			16'h0793;
		end
		32'h00009FFA: begin
				q			<=			16'h0240;
		end
		32'h00009FFC: begin
				q			<=			16'hE463;
		end
		32'h00009FFE: begin
				q			<=			16'h08C7;
		end
		32'h0000A000: begin
				q			<=			16'h0713;
		end
		32'h0000A002: begin
				q			<=			16'h0130;
		end
		32'h0000A004: begin
				q			<=			16'h7263;
		end
		32'h0000A006: begin
				q			<=			16'h02C7;
		end
		32'h0000A008: begin
				q			<=			16'h2703;
		end
		32'h0000A00A: begin
				q			<=			16'h0004;
		end
		32'h0000A00C: begin
				q			<=			16'hA423;
		end
		32'h0000A00E: begin
				q			<=			16'h00E4;
		end
		32'h0000A010: begin
				q			<=			16'h2703;
		end
		32'h0000A012: begin
				q			<=			16'h0044;
		end
		32'h0000A014: begin
				q			<=			16'hA623;
		end
		32'h0000A016: begin
				q			<=			16'h00E4;
		end
		32'h0000A018: begin
				q			<=			16'h0713;
		end
		32'h0000A01A: begin
				q			<=			16'h01B0;
		end
		32'h0000A01C: begin
				q			<=			16'h6663;
		end
		32'h0000A01E: begin
				q			<=			16'h02C7;
		end
		32'h0000A020: begin
				q			<=			16'h0413;
		end
		32'h0000A022: begin
				q			<=			16'h0084;
		end
		32'h0000A024: begin
				q			<=			16'h8513;
		end
		32'h0000A026: begin
				q			<=			16'h0104;
		end
		32'h0000A028: begin
				q			<=			16'h2783;
		end
		32'h0000A02A: begin
				q			<=			16'h0004;
		end
		32'h0000A02C: begin
				q			<=			16'h2023;
		end
		32'h0000A02E: begin
				q			<=			16'h00F5;
		end
		32'h0000A030: begin
				q			<=			16'h2783;
		end
		32'h0000A032: begin
				q			<=			16'h0044;
		end
		32'h0000A034: begin
				q			<=			16'h2223;
		end
		32'h0000A036: begin
				q			<=			16'h00F5;
		end
		32'h0000A038: begin
				q			<=			16'h2783;
		end
		32'h0000A03A: begin
				q			<=			16'h0084;
		end
		32'h0000A03C: begin
				q			<=			16'h2423;
		end
		32'h0000A03E: begin
				q			<=			16'h00F5;
		end
		32'h0000A040: begin
				q			<=			16'h0993;
		end
		32'h0000A042: begin
				q			<=			16'h000A;
		end
		32'h0000A044: begin
				q			<=			16'hF06F;
		end
		32'h0000A046: begin
				q			<=			16'hF49F;
		end
		32'h0000A048: begin
				q			<=			16'h2703;
		end
		32'h0000A04A: begin
				q			<=			16'h0084;
		end
		32'h0000A04C: begin
				q			<=			16'hA823;
		end
		32'h0000A04E: begin
				q			<=			16'h00E4;
		end
		32'h0000A050: begin
				q			<=			16'h2703;
		end
		32'h0000A052: begin
				q			<=			16'h00C4;
		end
		32'h0000A054: begin
				q			<=			16'hAA23;
		end
		32'h0000A056: begin
				q			<=			16'h00E4;
		end
		32'h0000A058: begin
				q			<=			16'h0863;
		end
		32'h0000A05A: begin
				q			<=			16'h00F6;
		end
		32'h0000A05C: begin
				q			<=			16'h0413;
		end
		32'h0000A05E: begin
				q			<=			16'h0104;
		end
		32'h0000A060: begin
				q			<=			16'h8513;
		end
		32'h0000A062: begin
				q			<=			16'h0184;
		end
		32'h0000A064: begin
				q			<=			16'hF06F;
		end
		32'h0000A066: begin
				q			<=			16'hFC5F;
		end
		32'h0000A068: begin
				q			<=			16'h2783;
		end
		32'h0000A06A: begin
				q			<=			16'h0104;
		end
		32'h0000A06C: begin
				q			<=			16'h8513;
		end
		32'h0000A06E: begin
				q			<=			16'h0204;
		end
		32'h0000A070: begin
				q			<=			16'h0413;
		end
		32'h0000A072: begin
				q			<=			16'h0184;
		end
		32'h0000A074: begin
				q			<=			16'hAC23;
		end
		32'h0000A076: begin
				q			<=			16'h00F4;
		end
		32'h0000A078: begin
				q			<=			16'h2783;
		end
		32'h0000A07A: begin
				q			<=			16'hFFC4;
		end
		32'h0000A07C: begin
				q			<=			16'hAE23;
		end
		32'h0000A07E: begin
				q			<=			16'h00F4;
		end
		32'h0000A080: begin
				q			<=			16'hF06F;
		end
		32'h0000A082: begin
				q			<=			16'hFA9F;
		end
		32'h0000A084: begin
				q			<=			16'h0593;
		end
		32'h0000A086: begin
				q			<=			16'h0004;
		end
		32'h0000A088: begin
				q			<=			16'hF0EF;
		end
		32'h0000A08A: begin
				q			<=			16'hB55F;
		end
		32'h0000A08C: begin
				q			<=			16'hF06F;
		end
		32'h0000A08E: begin
				q			<=			16'hFB5F;
		end
		32'h0000A090: begin
				q			<=			16'h8513;
		end
		32'h0000A092: begin
				q			<=			16'h000A;
		end
		32'h0000A094: begin
				q			<=			16'hD0EF;
		end
		32'h0000A096: begin
				q			<=			16'hB0CF;
		end
		32'h0000A098: begin
				q			<=			16'h0A13;
		end
		32'h0000A09A: begin
				q			<=			16'h0005;
		end
		32'h0000A09C: begin
				q			<=			16'h00E3;
		end
		32'h0000A09E: begin
				q			<=			16'hE205;
		end
		32'h0000A0A0: begin
				q			<=			16'h2783;
		end
		32'h0000A0A2: begin
				q			<=			16'hFFC4;
		end
		32'h0000A0A4: begin
				q			<=			16'h0713;
		end
		32'h0000A0A6: begin
				q			<=			16'hFF85;
		end
		32'h0000A0A8: begin
				q			<=			16'hF793;
		end
		32'h0000A0AA: begin
				q			<=			16'hFFE7;
		end
		32'h0000A0AC: begin
				q			<=			16'h87B3;
		end
		32'h0000A0AE: begin
				q			<=			16'h00FB;
		end
		32'h0000A0B0: begin
				q			<=			16'h9A63;
		end
		32'h0000A0B2: begin
				q			<=			16'h00E7;
		end
		32'h0000A0B4: begin
				q			<=			16'h2983;
		end
		32'h0000A0B6: begin
				q			<=			16'hFFC5;
		end
		32'h0000A0B8: begin
				q			<=			16'hF993;
		end
		32'h0000A0BA: begin
				q			<=			16'hFFC9;
		end
		32'h0000A0BC: begin
				q			<=			16'h89B3;
		end
		32'h0000A0BE: begin
				q			<=			16'h0129;
		end
		32'h0000A0C0: begin
				q			<=			16'hF06F;
		end
		32'h0000A0C2: begin
				q			<=			16'hCDDF;
		end
		32'h0000A0C4: begin
				q			<=			16'h0613;
		end
		32'h0000A0C6: begin
				q			<=			16'hFFC9;
		end
		32'h0000A0C8: begin
				q			<=			16'h0793;
		end
		32'h0000A0CA: begin
				q			<=			16'h0240;
		end
		32'h0000A0CC: begin
				q			<=			16'hE063;
		end
		32'h0000A0CE: begin
				q			<=			16'h0AC7;
		end
		32'h0000A0D0: begin
				q			<=			16'h0713;
		end
		32'h0000A0D2: begin
				q			<=			16'h0130;
		end
		32'h0000A0D4: begin
				q			<=			16'h7663;
		end
		32'h0000A0D6: begin
				q			<=			16'h08C7;
		end
		32'h0000A0D8: begin
				q			<=			16'h2703;
		end
		32'h0000A0DA: begin
				q			<=			16'h0004;
		end
		32'h0000A0DC: begin
				q			<=			16'h2023;
		end
		32'h0000A0DE: begin
				q			<=			16'h00E5;
		end
		32'h0000A0E0: begin
				q			<=			16'h2703;
		end
		32'h0000A0E2: begin
				q			<=			16'h0044;
		end
		32'h0000A0E4: begin
				q			<=			16'h2223;
		end
		32'h0000A0E6: begin
				q			<=			16'h00E5;
		end
		32'h0000A0E8: begin
				q			<=			16'h0713;
		end
		32'h0000A0EA: begin
				q			<=			16'h01B0;
		end
		32'h0000A0EC: begin
				q			<=			16'h6C63;
		end
		32'h0000A0EE: begin
				q			<=			16'h02C7;
		end
		32'h0000A0F0: begin
				q			<=			16'h0713;
		end
		32'h0000A0F2: begin
				q			<=			16'h0084;
		end
		32'h0000A0F4: begin
				q			<=			16'h0793;
		end
		32'h0000A0F6: begin
				q			<=			16'h0085;
		end
		32'h0000A0F8: begin
				q			<=			16'h2683;
		end
		32'h0000A0FA: begin
				q			<=			16'h0007;
		end
		32'h0000A0FC: begin
				q			<=			16'hA023;
		end
		32'h0000A0FE: begin
				q			<=			16'h00D7;
		end
		32'h0000A100: begin
				q			<=			16'h2683;
		end
		32'h0000A102: begin
				q			<=			16'h0047;
		end
		32'h0000A104: begin
				q			<=			16'hA223;
		end
		32'h0000A106: begin
				q			<=			16'h00D7;
		end
		32'h0000A108: begin
				q			<=			16'h2703;
		end
		32'h0000A10A: begin
				q			<=			16'h0087;
		end
		32'h0000A10C: begin
				q			<=			16'hA423;
		end
		32'h0000A10E: begin
				q			<=			16'h00E7;
		end
		32'h0000A110: begin
				q			<=			16'h0593;
		end
		32'h0000A112: begin
				q			<=			16'h0004;
		end
		32'h0000A114: begin
				q			<=			16'h8513;
		end
		32'h0000A116: begin
				q			<=			16'h000A;
		end
		32'h0000A118: begin
				q			<=			16'hB097;
		end
		32'h0000A11A: begin
				q			<=			16'hFFFF;
		end
		32'h0000A11C: begin
				q			<=			16'h80E7;
		end
		32'h0000A11E: begin
				q			<=			16'hE580;
		end
		32'h0000A120: begin
				q			<=			16'hF06F;
		end
		32'h0000A122: begin
				q			<=			16'hD9DF;
		end
		32'h0000A124: begin
				q			<=			16'h2703;
		end
		32'h0000A126: begin
				q			<=			16'h0084;
		end
		32'h0000A128: begin
				q			<=			16'h2423;
		end
		32'h0000A12A: begin
				q			<=			16'h00E5;
		end
		32'h0000A12C: begin
				q			<=			16'h2703;
		end
		32'h0000A12E: begin
				q			<=			16'h00C4;
		end
		32'h0000A130: begin
				q			<=			16'h2623;
		end
		32'h0000A132: begin
				q			<=			16'h00E5;
		end
		32'h0000A134: begin
				q			<=			16'h0863;
		end
		32'h0000A136: begin
				q			<=			16'h00F6;
		end
		32'h0000A138: begin
				q			<=			16'h0713;
		end
		32'h0000A13A: begin
				q			<=			16'h0104;
		end
		32'h0000A13C: begin
				q			<=			16'h0793;
		end
		32'h0000A13E: begin
				q			<=			16'h0105;
		end
		32'h0000A140: begin
				q			<=			16'hF06F;
		end
		32'h0000A142: begin
				q			<=			16'hFB9F;
		end
		32'h0000A144: begin
				q			<=			16'h2783;
		end
		32'h0000A146: begin
				q			<=			16'h0104;
		end
		32'h0000A148: begin
				q			<=			16'h0713;
		end
		32'h0000A14A: begin
				q			<=			16'h0184;
		end
		32'h0000A14C: begin
				q			<=			16'h2823;
		end
		32'h0000A14E: begin
				q			<=			16'h00F5;
		end
		32'h0000A150: begin
				q			<=			16'h2683;
		end
		32'h0000A152: begin
				q			<=			16'h0144;
		end
		32'h0000A154: begin
				q			<=			16'h0793;
		end
		32'h0000A156: begin
				q			<=			16'h0185;
		end
		32'h0000A158: begin
				q			<=			16'h2A23;
		end
		32'h0000A15A: begin
				q			<=			16'h00D5;
		end
		32'h0000A15C: begin
				q			<=			16'hF06F;
		end
		32'h0000A15E: begin
				q			<=			16'hF9DF;
		end
		32'h0000A160: begin
				q			<=			16'h0793;
		end
		32'h0000A162: begin
				q			<=			16'h0005;
		end
		32'h0000A164: begin
				q			<=			16'h0713;
		end
		32'h0000A166: begin
				q			<=			16'h0004;
		end
		32'h0000A168: begin
				q			<=			16'hF06F;
		end
		32'h0000A16A: begin
				q			<=			16'hF91F;
		end
		32'h0000A16C: begin
				q			<=			16'h0593;
		end
		32'h0000A16E: begin
				q			<=			16'h0004;
		end
		32'h0000A170: begin
				q			<=			16'hF0EF;
		end
		32'h0000A172: begin
				q			<=			16'hA6DF;
		end
		32'h0000A174: begin
				q			<=			16'hF06F;
		end
		32'h0000A176: begin
				q			<=			16'hF9DF;
		end
		32'h0000A178: begin
				q			<=			16'h0993;
		end
		32'h0000A17A: begin
				q			<=			16'h0009;
		end
		32'h0000A17C: begin
				q			<=			16'hF06F;
		end
		32'h0000A17E: begin
				q			<=			16'hC21F;
		end
		32'h0000A180: begin
				q			<=			16'hE9B3;
		end
		32'h0000A182: begin
				q			<=			16'h00E9;
		end
		32'h0000A184: begin
				q			<=			16'hA223;
		end
		32'h0000A186: begin
				q			<=			16'h013B;
		end
		32'h0000A188: begin
				q			<=			16'hA703;
		end
		32'h0000A18A: begin
				q			<=			16'h0047;
		end
		32'h0000A18C: begin
				q			<=			16'h6713;
		end
		32'h0000A18E: begin
				q			<=			16'h0017;
		end
		32'h0000A190: begin
				q			<=			16'hA223;
		end
		32'h0000A192: begin
				q			<=			16'h00E7;
		end
		32'h0000A194: begin
				q			<=			16'hF06F;
		end
		32'h0000A196: begin
				q			<=			16'hC51F;
		end
		32'h0000A198: begin
				q			<=			16'h0000;
		end
		32'h0000A19A: begin
				q			<=			16'h0000;
		end
		32'h0000A19C: begin
				q			<=			16'h0113;
		end
		32'h0000A19E: begin
				q			<=			16'hFF01;
		end
		32'h0000A1A0: begin
				q			<=			16'h2423;
		end
		32'h0000A1A2: begin
				q			<=			16'h0081;
		end
		32'h0000A1A4: begin
				q			<=			16'h8413;
		end
		32'h0000A1A6: begin
				q			<=			16'h0005;
		end
		32'h0000A1A8: begin
				q			<=			16'hA583;
		end
		32'h0000A1AA: begin
				q			<=			16'h0005;
		end
		32'h0000A1AC: begin
				q			<=			16'h2223;
		end
		32'h0000A1AE: begin
				q			<=			16'h0091;
		end
		32'h0000A1B0: begin
				q			<=			16'h2623;
		end
		32'h0000A1B2: begin
				q			<=			16'h0011;
		end
		32'h0000A1B4: begin
				q			<=			16'h0493;
		end
		32'h0000A1B6: begin
				q			<=			16'h0005;
		end
		32'h0000A1B8: begin
				q			<=			16'h8463;
		end
		32'h0000A1BA: begin
				q			<=			16'h0005;
		end
		32'h0000A1BC: begin
				q			<=			16'hF0EF;
		end
		32'h0000A1BE: begin
				q			<=			16'hFE1F;
		end
		32'h0000A1C0: begin
				q			<=			16'h0593;
		end
		32'h0000A1C2: begin
				q			<=			16'h0004;
		end
		32'h0000A1C4: begin
				q			<=			16'h2403;
		end
		32'h0000A1C6: begin
				q			<=			16'h0081;
		end
		32'h0000A1C8: begin
				q			<=			16'h2083;
		end
		32'h0000A1CA: begin
				q			<=			16'h00C1;
		end
		32'h0000A1CC: begin
				q			<=			16'h8513;
		end
		32'h0000A1CE: begin
				q			<=			16'h0004;
		end
		32'h0000A1D0: begin
				q			<=			16'h2483;
		end
		32'h0000A1D2: begin
				q			<=			16'h0041;
		end
		32'h0000A1D4: begin
				q			<=			16'h0113;
		end
		32'h0000A1D6: begin
				q			<=			16'h0101;
		end
		32'h0000A1D8: begin
				q			<=			16'hB317;
		end
		32'h0000A1DA: begin
				q			<=			16'hFFFF;
		end
		32'h0000A1DC: begin
				q			<=			16'h0067;
		end
		32'h0000A1DE: begin
				q			<=			16'hD983;
		end
		32'h0000A1E0: begin
				q			<=			16'h6797;
		end
		32'h0000A1E2: begin
				q			<=			16'h0000;
		end
		32'h0000A1E4: begin
				q			<=			16'h8793;
		end
		32'h0000A1E6: begin
				q			<=			16'h6F87;
		end
		32'h0000A1E8: begin
				q			<=			16'hA783;
		end
		32'h0000A1EA: begin
				q			<=			16'h0007;
		end
		32'h0000A1EC: begin
				q			<=			16'h8463;
		end
		32'h0000A1EE: begin
				q			<=			16'h10A7;
		end
		32'h0000A1F0: begin
				q			<=			16'h2783;
		end
		32'h0000A1F2: begin
				q			<=			16'h04C5;
		end
		32'h0000A1F4: begin
				q			<=			16'h0113;
		end
		32'h0000A1F6: begin
				q			<=			16'hFE01;
		end
		32'h0000A1F8: begin
				q			<=			16'h2C23;
		end
		32'h0000A1FA: begin
				q			<=			16'h0081;
		end
		32'h0000A1FC: begin
				q			<=			16'h2A23;
		end
		32'h0000A1FE: begin
				q			<=			16'h0091;
		end
		32'h0000A200: begin
				q			<=			16'h2823;
		end
		32'h0000A202: begin
				q			<=			16'h0121;
		end
		32'h0000A204: begin
				q			<=			16'h2E23;
		end
		32'h0000A206: begin
				q			<=			16'h0011;
		end
		32'h0000A208: begin
				q			<=			16'h2623;
		end
		32'h0000A20A: begin
				q			<=			16'h0131;
		end
		32'h0000A20C: begin
				q			<=			16'h0413;
		end
		32'h0000A20E: begin
				q			<=			16'h0005;
		end
		32'h0000A210: begin
				q			<=			16'h0493;
		end
		32'h0000A212: begin
				q			<=			16'h0000;
		end
		32'h0000A214: begin
				q			<=			16'h0913;
		end
		32'h0000A216: begin
				q			<=			16'h0800;
		end
		32'h0000A218: begin
				q			<=			16'h9463;
		end
		32'h0000A21A: begin
				q			<=			16'h0407;
		end
		32'h0000A21C: begin
				q			<=			16'h2583;
		end
		32'h0000A21E: begin
				q			<=			16'h0404;
		end
		32'h0000A220: begin
				q			<=			16'h8663;
		end
		32'h0000A222: begin
				q			<=			16'h0005;
		end
		32'h0000A224: begin
				q			<=			16'h0513;
		end
		32'h0000A226: begin
				q			<=			16'h0004;
		end
		32'h0000A228: begin
				q			<=			16'hA0EF;
		end
		32'h0000A22A: begin
				q			<=			16'hD49F;
		end
		32'h0000A22C: begin
				q			<=			16'h2583;
		end
		32'h0000A22E: begin
				q			<=			16'h1484;
		end
		32'h0000A230: begin
				q			<=			16'h8C63;
		end
		32'h0000A232: begin
				q			<=			16'h0405;
		end
		32'h0000A234: begin
				q			<=			16'h0493;
		end
		32'h0000A236: begin
				q			<=			16'h14C4;
		end
		32'h0000A238: begin
				q			<=			16'h8863;
		end
		32'h0000A23A: begin
				q			<=			16'h0495;
		end
		32'h0000A23C: begin
				q			<=			16'hA903;
		end
		32'h0000A23E: begin
				q			<=			16'h0005;
		end
		32'h0000A240: begin
				q			<=			16'h0513;
		end
		32'h0000A242: begin
				q			<=			16'h0004;
		end
		32'h0000A244: begin
				q			<=			16'hA0EF;
		end
		32'h0000A246: begin
				q			<=			16'hD2DF;
		end
		32'h0000A248: begin
				q			<=			16'h0593;
		end
		32'h0000A24A: begin
				q			<=			16'h0009;
		end
		32'h0000A24C: begin
				q			<=			16'hF06F;
		end
		32'h0000A24E: begin
				q			<=			16'hFEDF;
		end
		32'h0000A250: begin
				q			<=			16'h85B3;
		end
		32'h0000A252: begin
				q			<=			16'h0095;
		end
		32'h0000A254: begin
				q			<=			16'hA583;
		end
		32'h0000A256: begin
				q			<=			16'h0005;
		end
		32'h0000A258: begin
				q			<=			16'h9E63;
		end
		32'h0000A25A: begin
				q			<=			16'h0005;
		end
		32'h0000A25C: begin
				q			<=			16'h8493;
		end
		32'h0000A25E: begin
				q			<=			16'h0044;
		end
		32'h0000A260: begin
				q			<=			16'h2583;
		end
		32'h0000A262: begin
				q			<=			16'h04C4;
		end
		32'h0000A264: begin
				q			<=			16'h96E3;
		end
		32'h0000A266: begin
				q			<=			16'hFF24;
		end
		32'h0000A268: begin
				q			<=			16'h0513;
		end
		32'h0000A26A: begin
				q			<=			16'h0004;
		end
		32'h0000A26C: begin
				q			<=			16'hA0EF;
		end
		32'h0000A26E: begin
				q			<=			16'hD05F;
		end
		32'h0000A270: begin
				q			<=			16'hF06F;
		end
		32'h0000A272: begin
				q			<=			16'hFADF;
		end
		32'h0000A274: begin
				q			<=			16'hA983;
		end
		32'h0000A276: begin
				q			<=			16'h0005;
		end
		32'h0000A278: begin
				q			<=			16'h0513;
		end
		32'h0000A27A: begin
				q			<=			16'h0004;
		end
		32'h0000A27C: begin
				q			<=			16'hA0EF;
		end
		32'h0000A27E: begin
				q			<=			16'hCF5F;
		end
		32'h0000A280: begin
				q			<=			16'h8593;
		end
		32'h0000A282: begin
				q			<=			16'h0009;
		end
		32'h0000A284: begin
				q			<=			16'hF06F;
		end
		32'h0000A286: begin
				q			<=			16'hFD5F;
		end
		32'h0000A288: begin
				q			<=			16'h2583;
		end
		32'h0000A28A: begin
				q			<=			16'h0544;
		end
		32'h0000A28C: begin
				q			<=			16'h8663;
		end
		32'h0000A28E: begin
				q			<=			16'h0005;
		end
		32'h0000A290: begin
				q			<=			16'h0513;
		end
		32'h0000A292: begin
				q			<=			16'h0004;
		end
		32'h0000A294: begin
				q			<=			16'hA0EF;
		end
		32'h0000A296: begin
				q			<=			16'hCDDF;
		end
		32'h0000A298: begin
				q			<=			16'h2783;
		end
		32'h0000A29A: begin
				q			<=			16'h0384;
		end
		32'h0000A29C: begin
				q			<=			16'h8E63;
		end
		32'h0000A29E: begin
				q			<=			16'h0207;
		end
		32'h0000A2A0: begin
				q			<=			16'h2783;
		end
		32'h0000A2A2: begin
				q			<=			16'h03C4;
		end
		32'h0000A2A4: begin
				q			<=			16'h0513;
		end
		32'h0000A2A6: begin
				q			<=			16'h0004;
		end
		32'h0000A2A8: begin
				q			<=			16'h80E7;
		end
		32'h0000A2AA: begin
				q			<=			16'h0007;
		end
		32'h0000A2AC: begin
				q			<=			16'h2583;
		end
		32'h0000A2AE: begin
				q			<=			16'h2E04;
		end
		32'h0000A2B0: begin
				q			<=			16'h8463;
		end
		32'h0000A2B2: begin
				q			<=			16'h0205;
		end
		32'h0000A2B4: begin
				q			<=			16'h0513;
		end
		32'h0000A2B6: begin
				q			<=			16'h0004;
		end
		32'h0000A2B8: begin
				q			<=			16'h2403;
		end
		32'h0000A2BA: begin
				q			<=			16'h0181;
		end
		32'h0000A2BC: begin
				q			<=			16'h2083;
		end
		32'h0000A2BE: begin
				q			<=			16'h01C1;
		end
		32'h0000A2C0: begin
				q			<=			16'h2483;
		end
		32'h0000A2C2: begin
				q			<=			16'h0141;
		end
		32'h0000A2C4: begin
				q			<=			16'h2903;
		end
		32'h0000A2C6: begin
				q			<=			16'h0101;
		end
		32'h0000A2C8: begin
				q			<=			16'h2983;
		end
		32'h0000A2CA: begin
				q			<=			16'h00C1;
		end
		32'h0000A2CC: begin
				q			<=			16'h0113;
		end
		32'h0000A2CE: begin
				q			<=			16'h0201;
		end
		32'h0000A2D0: begin
				q			<=			16'h0317;
		end
		32'h0000A2D2: begin
				q			<=			16'h0000;
		end
		32'h0000A2D4: begin
				q			<=			16'h0067;
		end
		32'h0000A2D6: begin
				q			<=			16'hECC3;
		end
		32'h0000A2D8: begin
				q			<=			16'h2083;
		end
		32'h0000A2DA: begin
				q			<=			16'h01C1;
		end
		32'h0000A2DC: begin
				q			<=			16'h2403;
		end
		32'h0000A2DE: begin
				q			<=			16'h0181;
		end
		32'h0000A2E0: begin
				q			<=			16'h2483;
		end
		32'h0000A2E2: begin
				q			<=			16'h0141;
		end
		32'h0000A2E4: begin
				q			<=			16'h2903;
		end
		32'h0000A2E6: begin
				q			<=			16'h0101;
		end
		32'h0000A2E8: begin
				q			<=			16'h2983;
		end
		32'h0000A2EA: begin
				q			<=			16'h00C1;
		end
		32'h0000A2EC: begin
				q			<=			16'h0113;
		end
		32'h0000A2EE: begin
				q			<=			16'h0201;
		end
		32'h0000A2F0: begin
				q			<=			16'h8067;
		end
		32'h0000A2F2: begin
				q			<=			16'h0000;
		end
		32'h0000A2F4: begin
				q			<=			16'h8067;
		end
		32'h0000A2F6: begin
				q			<=			16'h0000;
		end
		32'h0000A2F8: begin
				q			<=			16'h0000;
		end
		32'h0000A2FA: begin
				q			<=			16'h0000;
		end
		32'h0000A2FC: begin
				q			<=			16'h6733;
		end
		32'h0000A2FE: begin
				q			<=			16'h00B5;
		end
		32'h0000A300: begin
				q			<=			16'h0393;
		end
		32'h0000A302: begin
				q			<=			16'hFFF0;
		end
		32'h0000A304: begin
				q			<=			16'h7713;
		end
		32'h0000A306: begin
				q			<=			16'h0037;
		end
		32'h0000A308: begin
				q			<=			16'h1063;
		end
		32'h0000A30A: begin
				q			<=			16'h1007;
		end
		32'h0000A30C: begin
				q			<=			16'h8E37;
		end
		32'h0000A30E: begin
				q			<=			16'h7F7F;
		end
		32'h0000A310: begin
				q			<=			16'h0E13;
		end
		32'h0000A312: begin
				q			<=			16'hF7FE;
		end
		32'h0000A314: begin
				q			<=			16'h2603;
		end
		32'h0000A316: begin
				q			<=			16'h0005;
		end
		32'h0000A318: begin
				q			<=			16'hA683;
		end
		32'h0000A31A: begin
				q			<=			16'h0005;
		end
		32'h0000A31C: begin
				q			<=			16'h72B3;
		end
		32'h0000A31E: begin
				q			<=			16'h01C6;
		end
		32'h0000A320: begin
				q			<=			16'h6333;
		end
		32'h0000A322: begin
				q			<=			16'h01C6;
		end
		32'h0000A324: begin
				q			<=			16'h82B3;
		end
		32'h0000A326: begin
				q			<=			16'h01C2;
		end
		32'h0000A328: begin
				q			<=			16'hE2B3;
		end
		32'h0000A32A: begin
				q			<=			16'h0062;
		end
		32'h0000A32C: begin
				q			<=			16'h9263;
		end
		32'h0000A32E: begin
				q			<=			16'h1072;
		end
		32'h0000A330: begin
				q			<=			16'h1663;
		end
		32'h0000A332: begin
				q			<=			16'h08D6;
		end
		32'h0000A334: begin
				q			<=			16'h2603;
		end
		32'h0000A336: begin
				q			<=			16'h0045;
		end
		32'h0000A338: begin
				q			<=			16'hA683;
		end
		32'h0000A33A: begin
				q			<=			16'h0045;
		end
		32'h0000A33C: begin
				q			<=			16'h72B3;
		end
		32'h0000A33E: begin
				q			<=			16'h01C6;
		end
		32'h0000A340: begin
				q			<=			16'h6333;
		end
		32'h0000A342: begin
				q			<=			16'h01C6;
		end
		32'h0000A344: begin
				q			<=			16'h82B3;
		end
		32'h0000A346: begin
				q			<=			16'h01C2;
		end
		32'h0000A348: begin
				q			<=			16'hE2B3;
		end
		32'h0000A34A: begin
				q			<=			16'h0062;
		end
		32'h0000A34C: begin
				q			<=			16'h9E63;
		end
		32'h0000A34E: begin
				q			<=			16'h0C72;
		end
		32'h0000A350: begin
				q			<=			16'h1663;
		end
		32'h0000A352: begin
				q			<=			16'h06D6;
		end
		32'h0000A354: begin
				q			<=			16'h2603;
		end
		32'h0000A356: begin
				q			<=			16'h0085;
		end
		32'h0000A358: begin
				q			<=			16'hA683;
		end
		32'h0000A35A: begin
				q			<=			16'h0085;
		end
		32'h0000A35C: begin
				q			<=			16'h72B3;
		end
		32'h0000A35E: begin
				q			<=			16'h01C6;
		end
		32'h0000A360: begin
				q			<=			16'h6333;
		end
		32'h0000A362: begin
				q			<=			16'h01C6;
		end
		32'h0000A364: begin
				q			<=			16'h82B3;
		end
		32'h0000A366: begin
				q			<=			16'h01C2;
		end
		32'h0000A368: begin
				q			<=			16'hE2B3;
		end
		32'h0000A36A: begin
				q			<=			16'h0062;
		end
		32'h0000A36C: begin
				q			<=			16'h9863;
		end
		32'h0000A36E: begin
				q			<=			16'h0C72;
		end
		32'h0000A370: begin
				q			<=			16'h1663;
		end
		32'h0000A372: begin
				q			<=			16'h04D6;
		end
		32'h0000A374: begin
				q			<=			16'h2603;
		end
		32'h0000A376: begin
				q			<=			16'h00C5;
		end
		32'h0000A378: begin
				q			<=			16'hA683;
		end
		32'h0000A37A: begin
				q			<=			16'h00C5;
		end
		32'h0000A37C: begin
				q			<=			16'h72B3;
		end
		32'h0000A37E: begin
				q			<=			16'h01C6;
		end
		32'h0000A380: begin
				q			<=			16'h6333;
		end
		32'h0000A382: begin
				q			<=			16'h01C6;
		end
		32'h0000A384: begin
				q			<=			16'h82B3;
		end
		32'h0000A386: begin
				q			<=			16'h01C2;
		end
		32'h0000A388: begin
				q			<=			16'hE2B3;
		end
		32'h0000A38A: begin
				q			<=			16'h0062;
		end
		32'h0000A38C: begin
				q			<=			16'h9263;
		end
		32'h0000A38E: begin
				q			<=			16'h0C72;
		end
		32'h0000A390: begin
				q			<=			16'h1663;
		end
		32'h0000A392: begin
				q			<=			16'h02D6;
		end
		32'h0000A394: begin
				q			<=			16'h2603;
		end
		32'h0000A396: begin
				q			<=			16'h0105;
		end
		32'h0000A398: begin
				q			<=			16'hA683;
		end
		32'h0000A39A: begin
				q			<=			16'h0105;
		end
		32'h0000A39C: begin
				q			<=			16'h72B3;
		end
		32'h0000A39E: begin
				q			<=			16'h01C6;
		end
		32'h0000A3A0: begin
				q			<=			16'h6333;
		end
		32'h0000A3A2: begin
				q			<=			16'h01C6;
		end
		32'h0000A3A4: begin
				q			<=			16'h82B3;
		end
		32'h0000A3A6: begin
				q			<=			16'h01C2;
		end
		32'h0000A3A8: begin
				q			<=			16'hE2B3;
		end
		32'h0000A3AA: begin
				q			<=			16'h0062;
		end
		32'h0000A3AC: begin
				q			<=			16'h9C63;
		end
		32'h0000A3AE: begin
				q			<=			16'h0A72;
		end
		32'h0000A3B0: begin
				q			<=			16'h0513;
		end
		32'h0000A3B2: begin
				q			<=			16'h0145;
		end
		32'h0000A3B4: begin
				q			<=			16'h8593;
		end
		32'h0000A3B6: begin
				q			<=			16'h0145;
		end
		32'h0000A3B8: begin
				q			<=			16'h0EE3;
		end
		32'h0000A3BA: begin
				q			<=			16'hF4D6;
		end
		32'h0000A3BC: begin
				q			<=			16'h1713;
		end
		32'h0000A3BE: begin
				q			<=			16'h0106;
		end
		32'h0000A3C0: begin
				q			<=			16'h9793;
		end
		32'h0000A3C2: begin
				q			<=			16'h0106;
		end
		32'h0000A3C4: begin
				q			<=			16'h1E63;
		end
		32'h0000A3C6: begin
				q			<=			16'h00F7;
		end
		32'h0000A3C8: begin
				q			<=			16'h5713;
		end
		32'h0000A3CA: begin
				q			<=			16'h0106;
		end
		32'h0000A3CC: begin
				q			<=			16'hD793;
		end
		32'h0000A3CE: begin
				q			<=			16'h0106;
		end
		32'h0000A3D0: begin
				q			<=			16'h0533;
		end
		32'h0000A3D2: begin
				q			<=			16'h40F7;
		end
		32'h0000A3D4: begin
				q			<=			16'h7593;
		end
		32'h0000A3D6: begin
				q			<=			16'h0FF5;
		end
		32'h0000A3D8: begin
				q			<=			16'h9063;
		end
		32'h0000A3DA: begin
				q			<=			16'h0205;
		end
		32'h0000A3DC: begin
				q			<=			16'h8067;
		end
		32'h0000A3DE: begin
				q			<=			16'h0000;
		end
		32'h0000A3E0: begin
				q			<=			16'h5713;
		end
		32'h0000A3E2: begin
				q			<=			16'h0107;
		end
		32'h0000A3E4: begin
				q			<=			16'hD793;
		end
		32'h0000A3E6: begin
				q			<=			16'h0107;
		end
		32'h0000A3E8: begin
				q			<=			16'h0533;
		end
		32'h0000A3EA: begin
				q			<=			16'h40F7;
		end
		32'h0000A3EC: begin
				q			<=			16'h7593;
		end
		32'h0000A3EE: begin
				q			<=			16'h0FF5;
		end
		32'h0000A3F0: begin
				q			<=			16'h9463;
		end
		32'h0000A3F2: begin
				q			<=			16'h0005;
		end
		32'h0000A3F4: begin
				q			<=			16'h8067;
		end
		32'h0000A3F6: begin
				q			<=			16'h0000;
		end
		32'h0000A3F8: begin
				q			<=			16'h7713;
		end
		32'h0000A3FA: begin
				q			<=			16'h0FF7;
		end
		32'h0000A3FC: begin
				q			<=			16'hF793;
		end
		32'h0000A3FE: begin
				q			<=			16'h0FF7;
		end
		32'h0000A400: begin
				q			<=			16'h0533;
		end
		32'h0000A402: begin
				q			<=			16'h40F7;
		end
		32'h0000A404: begin
				q			<=			16'h8067;
		end
		32'h0000A406: begin
				q			<=			16'h0000;
		end
		32'h0000A408: begin
				q			<=			16'h4603;
		end
		32'h0000A40A: begin
				q			<=			16'h0005;
		end
		32'h0000A40C: begin
				q			<=			16'hC683;
		end
		32'h0000A40E: begin
				q			<=			16'h0005;
		end
		32'h0000A410: begin
				q			<=			16'h0513;
		end
		32'h0000A412: begin
				q			<=			16'h0015;
		end
		32'h0000A414: begin
				q			<=			16'h8593;
		end
		32'h0000A416: begin
				q			<=			16'h0015;
		end
		32'h0000A418: begin
				q			<=			16'h1463;
		end
		32'h0000A41A: begin
				q			<=			16'h00D6;
		end
		32'h0000A41C: begin
				q			<=			16'h16E3;
		end
		32'h0000A41E: begin
				q			<=			16'hFE06;
		end
		32'h0000A420: begin
				q			<=			16'h0533;
		end
		32'h0000A422: begin
				q			<=			16'h40D6;
		end
		32'h0000A424: begin
				q			<=			16'h8067;
		end
		32'h0000A426: begin
				q			<=			16'h0000;
		end
		32'h0000A428: begin
				q			<=			16'h0513;
		end
		32'h0000A42A: begin
				q			<=			16'h0045;
		end
		32'h0000A42C: begin
				q			<=			16'h8593;
		end
		32'h0000A42E: begin
				q			<=			16'h0045;
		end
		32'h0000A430: begin
				q			<=			16'h1CE3;
		end
		32'h0000A432: begin
				q			<=			16'hFCD6;
		end
		32'h0000A434: begin
				q			<=			16'h0513;
		end
		32'h0000A436: begin
				q			<=			16'h0000;
		end
		32'h0000A438: begin
				q			<=			16'h8067;
		end
		32'h0000A43A: begin
				q			<=			16'h0000;
		end
		32'h0000A43C: begin
				q			<=			16'h0513;
		end
		32'h0000A43E: begin
				q			<=			16'h0085;
		end
		32'h0000A440: begin
				q			<=			16'h8593;
		end
		32'h0000A442: begin
				q			<=			16'h0085;
		end
		32'h0000A444: begin
				q			<=			16'h12E3;
		end
		32'h0000A446: begin
				q			<=			16'hFCD6;
		end
		32'h0000A448: begin
				q			<=			16'h0513;
		end
		32'h0000A44A: begin
				q			<=			16'h0000;
		end
		32'h0000A44C: begin
				q			<=			16'h8067;
		end
		32'h0000A44E: begin
				q			<=			16'h0000;
		end
		32'h0000A450: begin
				q			<=			16'h0513;
		end
		32'h0000A452: begin
				q			<=			16'h00C5;
		end
		32'h0000A454: begin
				q			<=			16'h8593;
		end
		32'h0000A456: begin
				q			<=			16'h00C5;
		end
		32'h0000A458: begin
				q			<=			16'h18E3;
		end
		32'h0000A45A: begin
				q			<=			16'hFAD6;
		end
		32'h0000A45C: begin
				q			<=			16'h0513;
		end
		32'h0000A45E: begin
				q			<=			16'h0000;
		end
		32'h0000A460: begin
				q			<=			16'h8067;
		end
		32'h0000A462: begin
				q			<=			16'h0000;
		end
		32'h0000A464: begin
				q			<=			16'h0513;
		end
		32'h0000A466: begin
				q			<=			16'h0105;
		end
		32'h0000A468: begin
				q			<=			16'h8593;
		end
		32'h0000A46A: begin
				q			<=			16'h0105;
		end
		32'h0000A46C: begin
				q			<=			16'h1EE3;
		end
		32'h0000A46E: begin
				q			<=			16'hF8D6;
		end
		32'h0000A470: begin
				q			<=			16'h0513;
		end
		32'h0000A472: begin
				q			<=			16'h0000;
		end
		32'h0000A474: begin
				q			<=			16'h8067;
		end
		32'h0000A476: begin
				q			<=			16'h0000;
		end
		32'h0000A478: begin
				q			<=			16'h6797;
		end
		32'h0000A47A: begin
				q			<=			16'h0000;
		end
		32'h0000A47C: begin
				q			<=			16'h8793;
		end
		32'h0000A47E: begin
				q			<=			16'h4607;
		end
		32'h0000A480: begin
				q			<=			16'hA783;
		end
		32'h0000A482: begin
				q			<=			16'h0007;
		end
		32'h0000A484: begin
				q			<=			16'hA783;
		end
		32'h0000A486: begin
				q			<=			16'h0347;
		end
		32'h0000A488: begin
				q			<=			16'h9663;
		end
		32'h0000A48A: begin
				q			<=			16'h0007;
		end
		32'h0000A48C: begin
				q			<=			16'h6797;
		end
		32'h0000A48E: begin
				q			<=			16'h0000;
		end
		32'h0000A490: begin
				q			<=			16'h8793;
		end
		32'h0000A492: begin
				q			<=			16'h2DC7;
		end
		32'h0000A494: begin
				q			<=			16'hA303;
		end
		32'h0000A496: begin
				q			<=			16'h0E07;
		end
		32'h0000A498: begin
				q			<=			16'h0067;
		end
		32'h0000A49A: begin
				q			<=			16'h0003;
		end
		32'h0000A49C: begin
				q			<=			16'h8463;
		end
		32'h0000A49E: begin
				q			<=			16'h0205;
		end
		32'h0000A4A0: begin
				q			<=			16'h0793;
		end
		32'h0000A4A2: begin
				q			<=			16'h0FF0;
		end
		32'h0000A4A4: begin
				q			<=			16'hFA63;
		end
		32'h0000A4A6: begin
				q			<=			16'h00C7;
		end
		32'h0000A4A8: begin
				q			<=			16'h0793;
		end
		32'h0000A4AA: begin
				q			<=			16'h08A0;
		end
		32'h0000A4AC: begin
				q			<=			16'h2023;
		end
		32'h0000A4AE: begin
				q			<=			16'h00F5;
		end
		32'h0000A4B0: begin
				q			<=			16'h0513;
		end
		32'h0000A4B2: begin
				q			<=			16'hFFF0;
		end
		32'h0000A4B4: begin
				q			<=			16'h8067;
		end
		32'h0000A4B6: begin
				q			<=			16'h0000;
		end
		32'h0000A4B8: begin
				q			<=			16'h8023;
		end
		32'h0000A4BA: begin
				q			<=			16'h00C5;
		end
		32'h0000A4BC: begin
				q			<=			16'h0513;
		end
		32'h0000A4BE: begin
				q			<=			16'h0010;
		end
		32'h0000A4C0: begin
				q			<=			16'h8067;
		end
		32'h0000A4C2: begin
				q			<=			16'h0000;
		end
		32'h0000A4C4: begin
				q			<=			16'h0513;
		end
		32'h0000A4C6: begin
				q			<=			16'h0000;
		end
		32'h0000A4C8: begin
				q			<=			16'h8067;
		end
		32'h0000A4CA: begin
				q			<=			16'h0000;
		end
		32'h0000A4CC: begin
				q			<=			16'h0000;
		end
		32'h0000A4CE: begin
				q			<=			16'h0000;
		end
		32'h0000A4D0: begin
				q			<=			16'hA783;
		end
		32'h0000A4D2: begin
				q			<=			16'h0005;
		end
		32'h0000A4D4: begin
				q			<=			16'h1023;
		end
		32'h0000A4D6: begin
				q			<=			16'h00F5;
		end
		32'h0000A4D8: begin
				q			<=			16'hA783;
		end
		32'h0000A4DA: begin
				q			<=			16'h0085;
		end
		32'h0000A4DC: begin
				q			<=			16'h1123;
		end
		32'h0000A4DE: begin
				q			<=			16'h00F5;
		end
		32'h0000A4E0: begin
				q			<=			16'hA783;
		end
		32'h0000A4E2: begin
				q			<=			16'h0105;
		end
		32'h0000A4E4: begin
				q			<=			16'h2223;
		end
		32'h0000A4E6: begin
				q			<=			16'h00F5;
		end
		32'h0000A4E8: begin
				q			<=			16'hA783;
		end
		32'h0000A4EA: begin
				q			<=			16'h0145;
		end
		32'h0000A4EC: begin
				q			<=			16'h1423;
		end
		32'h0000A4EE: begin
				q			<=			16'h00F5;
		end
		32'h0000A4F0: begin
				q			<=			16'hA783;
		end
		32'h0000A4F2: begin
				q			<=			16'h0185;
		end
		32'h0000A4F4: begin
				q			<=			16'h1523;
		end
		32'h0000A4F6: begin
				q			<=			16'h00F5;
		end
		32'h0000A4F8: begin
				q			<=			16'hA783;
		end
		32'h0000A4FA: begin
				q			<=			16'h01C5;
		end
		32'h0000A4FC: begin
				q			<=			16'h1623;
		end
		32'h0000A4FE: begin
				q			<=			16'h00F5;
		end
		32'h0000A500: begin
				q			<=			16'hA783;
		end
		32'h0000A502: begin
				q			<=			16'h0205;
		end
		32'h0000A504: begin
				q			<=			16'h1723;
		end
		32'h0000A506: begin
				q			<=			16'h00F5;
		end
		32'h0000A508: begin
				q			<=			16'hA783;
		end
		32'h0000A50A: begin
				q			<=			16'h0305;
		end
		32'h0000A50C: begin
				q			<=			16'h2823;
		end
		32'h0000A50E: begin
				q			<=			16'h00F5;
		end
		32'h0000A510: begin
				q			<=			16'hA783;
		end
		32'h0000A512: begin
				q			<=			16'h0405;
		end
		32'h0000A514: begin
				q			<=			16'h2823;
		end
		32'h0000A516: begin
				q			<=			16'h02F5;
		end
		32'h0000A518: begin
				q			<=			16'hA783;
		end
		32'h0000A51A: begin
				q			<=			16'h0385;
		end
		32'h0000A51C: begin
				q			<=			16'h2623;
		end
		32'h0000A51E: begin
				q			<=			16'h02F5;
		end
		32'h0000A520: begin
				q			<=			16'hA783;
		end
		32'h0000A522: begin
				q			<=			16'h0485;
		end
		32'h0000A524: begin
				q			<=			16'h2A23;
		end
		32'h0000A526: begin
				q			<=			16'h00F5;
		end
		32'h0000A528: begin
				q			<=			16'hA783;
		end
		32'h0000A52A: begin
				q			<=			16'h0505;
		end
		32'h0000A52C: begin
				q			<=			16'h2E23;
		end
		32'h0000A52E: begin
				q			<=			16'h00F5;
		end
		32'h0000A530: begin
				q			<=			16'hA783;
		end
		32'h0000A532: begin
				q			<=			16'h0585;
		end
		32'h0000A534: begin
				q			<=			16'h2223;
		end
		32'h0000A536: begin
				q			<=			16'h02F5;
		end
		32'h0000A538: begin
				q			<=			16'h8067;
		end
		32'h0000A53A: begin
				q			<=			16'h0000;
		end
		32'h0000A53C: begin
				q			<=			16'h0113;
		end
		32'h0000A53E: begin
				q			<=			16'hFF01;
		end
		32'h0000A540: begin
				q			<=			16'h2423;
		end
		32'h0000A542: begin
				q			<=			16'h0081;
		end
		32'h0000A544: begin
				q			<=			16'h2623;
		end
		32'h0000A546: begin
				q			<=			16'h0011;
		end
		32'h0000A548: begin
				q			<=			16'h0413;
		end
		32'h0000A54A: begin
				q			<=			16'h0005;
		end
		32'h0000A54C: begin
				q			<=			16'h0097;
		end
		32'h0000A54E: begin
				q			<=			16'h0000;
		end
		32'h0000A550: begin
				q			<=			16'h80E7;
		end
		32'h0000A552: begin
				q			<=			16'h54C0;
		end
		32'h0000A554: begin
				q			<=			16'h07B3;
		end
		32'h0000A556: begin
				q			<=			16'h4080;
		end
		32'h0000A558: begin
				q			<=			16'h2083;
		end
		32'h0000A55A: begin
				q			<=			16'h00C1;
		end
		32'h0000A55C: begin
				q			<=			16'h2403;
		end
		32'h0000A55E: begin
				q			<=			16'h0081;
		end
		32'h0000A560: begin
				q			<=			16'h2023;
		end
		32'h0000A562: begin
				q			<=			16'h00F5;
		end
		32'h0000A564: begin
				q			<=			16'h0513;
		end
		32'h0000A566: begin
				q			<=			16'hFFF0;
		end
		32'h0000A568: begin
				q			<=			16'h0113;
		end
		32'h0000A56A: begin
				q			<=			16'h0101;
		end
		32'h0000A56C: begin
				q			<=			16'h8067;
		end
		32'h0000A56E: begin
				q			<=			16'h0000;
		end
		32'h0000A570: begin
				q			<=			16'h0893;
		end
		32'h0000A572: begin
				q			<=			16'h0005;
		end
		32'h0000A574: begin
				q			<=			16'h8513;
		end
		32'h0000A576: begin
				q			<=			16'h0005;
		end
		32'h0000A578: begin
				q			<=			16'h0593;
		end
		32'h0000A57A: begin
				q			<=			16'h0006;
		end
		32'h0000A57C: begin
				q			<=			16'h8613;
		end
		32'h0000A57E: begin
				q			<=			16'h0006;
		end
		32'h0000A580: begin
				q			<=			16'h0693;
		end
		32'h0000A582: begin
				q			<=			16'h0007;
		end
		32'h0000A584: begin
				q			<=			16'h0073;
		end
		32'h0000A586: begin
				q			<=			16'h0000;
		end
		32'h0000A588: begin
				q			<=			16'h5663;
		end
		32'h0000A58A: begin
				q			<=			16'h0005;
		end
		32'h0000A58C: begin
				q			<=			16'h0317;
		end
		32'h0000A58E: begin
				q			<=			16'h0000;
		end
		32'h0000A590: begin
				q			<=			16'h0067;
		end
		32'h0000A592: begin
				q			<=			16'hFB03;
		end
		32'h0000A594: begin
				q			<=			16'h8067;
		end
		32'h0000A596: begin
				q			<=			16'h0000;
		end
		32'h0000A598: begin
				q			<=			16'h0693;
		end
		32'h0000A59A: begin
				q			<=			16'h0006;
		end
		32'h0000A59C: begin
				q			<=			16'h0713;
		end
		32'h0000A59E: begin
				q			<=			16'h0000;
		end
		32'h0000A5A0: begin
				q			<=			16'h8613;
		end
		32'h0000A5A2: begin
				q			<=			16'h0005;
		end
		32'h0000A5A4: begin
				q			<=			16'h0593;
		end
		32'h0000A5A6: begin
				q			<=			16'h0005;
		end
		32'h0000A5A8: begin
				q			<=			16'h0513;
		end
		32'h0000A5AA: begin
				q			<=			16'h4000;
		end
		32'h0000A5AC: begin
				q			<=			16'h0317;
		end
		32'h0000A5AE: begin
				q			<=			16'h0000;
		end
		32'h0000A5B0: begin
				q			<=			16'h0067;
		end
		32'h0000A5B2: begin
				q			<=			16'hFC43;
		end
		32'h0000A5B4: begin
				q			<=			16'h8713;
		end
		32'h0000A5B6: begin
				q			<=			16'h0006;
		end
		32'h0000A5B8: begin
				q			<=			16'h0693;
		end
		32'h0000A5BA: begin
				q			<=			16'h0006;
		end
		32'h0000A5BC: begin
				q			<=			16'h8613;
		end
		32'h0000A5BE: begin
				q			<=			16'h0005;
		end
		32'h0000A5C0: begin
				q			<=			16'h0593;
		end
		32'h0000A5C2: begin
				q			<=			16'h0005;
		end
		32'h0000A5C4: begin
				q			<=			16'h0513;
		end
		32'h0000A5C6: begin
				q			<=			16'h0380;
		end
		32'h0000A5C8: begin
				q			<=			16'hF06F;
		end
		32'h0000A5CA: begin
				q			<=			16'hFA9F;
		end
		32'h0000A5CC: begin
				q			<=			16'h0693;
		end
		32'h0000A5CE: begin
				q			<=			16'h0006;
		end
		32'h0000A5D0: begin
				q			<=			16'h0713;
		end
		32'h0000A5D2: begin
				q			<=			16'h0000;
		end
		32'h0000A5D4: begin
				q			<=			16'h8613;
		end
		32'h0000A5D6: begin
				q			<=			16'h0005;
		end
		32'h0000A5D8: begin
				q			<=			16'h0593;
		end
		32'h0000A5DA: begin
				q			<=			16'h0005;
		end
		32'h0000A5DC: begin
				q			<=			16'h0513;
		end
		32'h0000A5DE: begin
				q			<=			16'h03E0;
		end
		32'h0000A5E0: begin
				q			<=			16'h0317;
		end
		32'h0000A5E2: begin
				q			<=			16'h0000;
		end
		32'h0000A5E4: begin
				q			<=			16'h0067;
		end
		32'h0000A5E6: begin
				q			<=			16'hF903;
		end
		32'h0000A5E8: begin
				q			<=			16'h0693;
		end
		32'h0000A5EA: begin
				q			<=			16'h0006;
		end
		32'h0000A5EC: begin
				q			<=			16'h0713;
		end
		32'h0000A5EE: begin
				q			<=			16'h0000;
		end
		32'h0000A5F0: begin
				q			<=			16'h8613;
		end
		32'h0000A5F2: begin
				q			<=			16'h0005;
		end
		32'h0000A5F4: begin
				q			<=			16'h0593;
		end
		32'h0000A5F6: begin
				q			<=			16'h0005;
		end
		32'h0000A5F8: begin
				q			<=			16'h0513;
		end
		32'h0000A5FA: begin
				q			<=			16'h03F0;
		end
		32'h0000A5FC: begin
				q			<=			16'hF06F;
		end
		32'h0000A5FE: begin
				q			<=			16'hF75F;
		end
		32'h0000A600: begin
				q			<=			16'h0693;
		end
		32'h0000A602: begin
				q			<=			16'h0006;
		end
		32'h0000A604: begin
				q			<=			16'h0713;
		end
		32'h0000A606: begin
				q			<=			16'h0000;
		end
		32'h0000A608: begin
				q			<=			16'h8613;
		end
		32'h0000A60A: begin
				q			<=			16'h0005;
		end
		32'h0000A60C: begin
				q			<=			16'h0593;
		end
		32'h0000A60E: begin
				q			<=			16'h0005;
		end
		32'h0000A610: begin
				q			<=			16'h0513;
		end
		32'h0000A612: begin
				q			<=			16'h0400;
		end
		32'h0000A614: begin
				q			<=			16'h0317;
		end
		32'h0000A616: begin
				q			<=			16'h0000;
		end
		32'h0000A618: begin
				q			<=			16'h0067;
		end
		32'h0000A61A: begin
				q			<=			16'hF5C3;
		end
		32'h0000A61C: begin
				q			<=			16'h0113;
		end
		32'h0000A61E: begin
				q			<=			16'hF801;
		end
		32'h0000A620: begin
				q			<=			16'h2A23;
		end
		32'h0000A622: begin
				q			<=			16'h0691;
		end
		32'h0000A624: begin
				q			<=			16'h0613;
		end
		32'h0000A626: begin
				q			<=			16'h0081;
		end
		32'h0000A628: begin
				q			<=			16'h8493;
		end
		32'h0000A62A: begin
				q			<=			16'h0005;
		end
		32'h0000A62C: begin
				q			<=			16'h0713;
		end
		32'h0000A62E: begin
				q			<=			16'h0000;
		end
		32'h0000A630: begin
				q			<=			16'h0593;
		end
		32'h0000A632: begin
				q			<=			16'h0005;
		end
		32'h0000A634: begin
				q			<=			16'h0693;
		end
		32'h0000A636: begin
				q			<=			16'h0000;
		end
		32'h0000A638: begin
				q			<=			16'h0513;
		end
		32'h0000A63A: begin
				q			<=			16'h0500;
		end
		32'h0000A63C: begin
				q			<=			16'h2E23;
		end
		32'h0000A63E: begin
				q			<=			16'h0611;
		end
		32'h0000A640: begin
				q			<=			16'h2C23;
		end
		32'h0000A642: begin
				q			<=			16'h0681;
		end
		32'h0000A644: begin
				q			<=			16'hF0EF;
		end
		32'h0000A646: begin
				q			<=			16'hF2DF;
		end
		32'h0000A648: begin
				q			<=			16'h0413;
		end
		32'h0000A64A: begin
				q			<=			16'h0005;
		end
		32'h0000A64C: begin
				q			<=			16'h0593;
		end
		32'h0000A64E: begin
				q			<=			16'h0081;
		end
		32'h0000A650: begin
				q			<=			16'h8513;
		end
		32'h0000A652: begin
				q			<=			16'h0004;
		end
		32'h0000A654: begin
				q			<=			16'hF0EF;
		end
		32'h0000A656: begin
				q			<=			16'hE7DF;
		end
		32'h0000A658: begin
				q			<=			16'h0513;
		end
		32'h0000A65A: begin
				q			<=			16'h0004;
		end
		32'h0000A65C: begin
				q			<=			16'h2083;
		end
		32'h0000A65E: begin
				q			<=			16'h07C1;
		end
		32'h0000A660: begin
				q			<=			16'h2403;
		end
		32'h0000A662: begin
				q			<=			16'h0781;
		end
		32'h0000A664: begin
				q			<=			16'h2483;
		end
		32'h0000A666: begin
				q			<=			16'h0741;
		end
		32'h0000A668: begin
				q			<=			16'h0113;
		end
		32'h0000A66A: begin
				q			<=			16'h0801;
		end
		32'h0000A66C: begin
				q			<=			16'h8067;
		end
		32'h0000A66E: begin
				q			<=			16'h0000;
		end
		32'h0000A670: begin
				q			<=			16'h0113;
		end
		32'h0000A672: begin
				q			<=			16'hF801;
		end
		32'h0000A674: begin
				q			<=			16'h2A23;
		end
		32'h0000A676: begin
				q			<=			16'h0691;
		end
		32'h0000A678: begin
				q			<=			16'h0613;
		end
		32'h0000A67A: begin
				q			<=			16'h0081;
		end
		32'h0000A67C: begin
				q			<=			16'h8493;
		end
		32'h0000A67E: begin
				q			<=			16'h0005;
		end
		32'h0000A680: begin
				q			<=			16'h0713;
		end
		32'h0000A682: begin
				q			<=			16'h0000;
		end
		32'h0000A684: begin
				q			<=			16'h0593;
		end
		32'h0000A686: begin
				q			<=			16'h0005;
		end
		32'h0000A688: begin
				q			<=			16'h0693;
		end
		32'h0000A68A: begin
				q			<=			16'h0000;
		end
		32'h0000A68C: begin
				q			<=			16'h0513;
		end
		32'h0000A68E: begin
				q			<=			16'h40E0;
		end
		32'h0000A690: begin
				q			<=			16'h2E23;
		end
		32'h0000A692: begin
				q			<=			16'h0611;
		end
		32'h0000A694: begin
				q			<=			16'h2C23;
		end
		32'h0000A696: begin
				q			<=			16'h0681;
		end
		32'h0000A698: begin
				q			<=			16'h0097;
		end
		32'h0000A69A: begin
				q			<=			16'h0000;
		end
		32'h0000A69C: begin
				q			<=			16'h80E7;
		end
		32'h0000A69E: begin
				q			<=			16'hED80;
		end
		32'h0000A6A0: begin
				q			<=			16'h0413;
		end
		32'h0000A6A2: begin
				q			<=			16'h0005;
		end
		32'h0000A6A4: begin
				q			<=			16'h0593;
		end
		32'h0000A6A6: begin
				q			<=			16'h0081;
		end
		32'h0000A6A8: begin
				q			<=			16'h8513;
		end
		32'h0000A6AA: begin
				q			<=			16'h0004;
		end
		32'h0000A6AC: begin
				q			<=			16'h0097;
		end
		32'h0000A6AE: begin
				q			<=			16'h0000;
		end
		32'h0000A6B0: begin
				q			<=			16'h80E7;
		end
		32'h0000A6B2: begin
				q			<=			16'hE240;
		end
		32'h0000A6B4: begin
				q			<=			16'h0513;
		end
		32'h0000A6B6: begin
				q			<=			16'h0004;
		end
		32'h0000A6B8: begin
				q			<=			16'h2083;
		end
		32'h0000A6BA: begin
				q			<=			16'h07C1;
		end
		32'h0000A6BC: begin
				q			<=			16'h2403;
		end
		32'h0000A6BE: begin
				q			<=			16'h0781;
		end
		32'h0000A6C0: begin
				q			<=			16'h2483;
		end
		32'h0000A6C2: begin
				q			<=			16'h0741;
		end
		32'h0000A6C4: begin
				q			<=			16'h0113;
		end
		32'h0000A6C6: begin
				q			<=			16'h0801;
		end
		32'h0000A6C8: begin
				q			<=			16'h8067;
		end
		32'h0000A6CA: begin
				q			<=			16'h0000;
		end
		32'h0000A6CC: begin
				q			<=			16'h0113;
		end
		32'h0000A6CE: begin
				q			<=			16'hF801;
		end
		32'h0000A6D0: begin
				q			<=			16'h2A23;
		end
		32'h0000A6D2: begin
				q			<=			16'h0691;
		end
		32'h0000A6D4: begin
				q			<=			16'h0613;
		end
		32'h0000A6D6: begin
				q			<=			16'h0081;
		end
		32'h0000A6D8: begin
				q			<=			16'h8493;
		end
		32'h0000A6DA: begin
				q			<=			16'h0005;
		end
		32'h0000A6DC: begin
				q			<=			16'h0713;
		end
		32'h0000A6DE: begin
				q			<=			16'h0000;
		end
		32'h0000A6E0: begin
				q			<=			16'h0593;
		end
		32'h0000A6E2: begin
				q			<=			16'h0005;
		end
		32'h0000A6E4: begin
				q			<=			16'h0693;
		end
		32'h0000A6E6: begin
				q			<=			16'h0000;
		end
		32'h0000A6E8: begin
				q			<=			16'h0513;
		end
		32'h0000A6EA: begin
				q			<=			16'h40F0;
		end
		32'h0000A6EC: begin
				q			<=			16'h2E23;
		end
		32'h0000A6EE: begin
				q			<=			16'h0611;
		end
		32'h0000A6F0: begin
				q			<=			16'h2C23;
		end
		32'h0000A6F2: begin
				q			<=			16'h0681;
		end
		32'h0000A6F4: begin
				q			<=			16'hF0EF;
		end
		32'h0000A6F6: begin
				q			<=			16'hE7DF;
		end
		32'h0000A6F8: begin
				q			<=			16'h0413;
		end
		32'h0000A6FA: begin
				q			<=			16'h0005;
		end
		32'h0000A6FC: begin
				q			<=			16'h0593;
		end
		32'h0000A6FE: begin
				q			<=			16'h0081;
		end
		32'h0000A700: begin
				q			<=			16'h8513;
		end
		32'h0000A702: begin
				q			<=			16'h0004;
		end
		32'h0000A704: begin
				q			<=			16'hF0EF;
		end
		32'h0000A706: begin
				q			<=			16'hDCDF;
		end
		32'h0000A708: begin
				q			<=			16'h0513;
		end
		32'h0000A70A: begin
				q			<=			16'h0004;
		end
		32'h0000A70C: begin
				q			<=			16'h2083;
		end
		32'h0000A70E: begin
				q			<=			16'h07C1;
		end
		32'h0000A710: begin
				q			<=			16'h2403;
		end
		32'h0000A712: begin
				q			<=			16'h0781;
		end
		32'h0000A714: begin
				q			<=			16'h2483;
		end
		32'h0000A716: begin
				q			<=			16'h0741;
		end
		32'h0000A718: begin
				q			<=			16'h0113;
		end
		32'h0000A71A: begin
				q			<=			16'h0801;
		end
		32'h0000A71C: begin
				q			<=			16'h8067;
		end
		32'h0000A71E: begin
				q			<=			16'h0000;
		end
		32'h0000A720: begin
				q			<=			16'h0113;
		end
		32'h0000A722: begin
				q			<=			16'hF801;
		end
		32'h0000A724: begin
				q			<=			16'h2A23;
		end
		32'h0000A726: begin
				q			<=			16'h0691;
		end
		32'h0000A728: begin
				q			<=			16'h8713;
		end
		32'h0000A72A: begin
				q			<=			16'h0006;
		end
		32'h0000A72C: begin
				q			<=			16'h0493;
		end
		32'h0000A72E: begin
				q			<=			16'h0006;
		end
		32'h0000A730: begin
				q			<=			16'h0693;
		end
		32'h0000A732: begin
				q			<=			16'h0081;
		end
		32'h0000A734: begin
				q			<=			16'h8613;
		end
		32'h0000A736: begin
				q			<=			16'h0005;
		end
		32'h0000A738: begin
				q			<=			16'h0593;
		end
		32'h0000A73A: begin
				q			<=			16'h0005;
		end
		32'h0000A73C: begin
				q			<=			16'h0513;
		end
		32'h0000A73E: begin
				q			<=			16'h04F0;
		end
		32'h0000A740: begin
				q			<=			16'h2E23;
		end
		32'h0000A742: begin
				q			<=			16'h0611;
		end
		32'h0000A744: begin
				q			<=			16'h2C23;
		end
		32'h0000A746: begin
				q			<=			16'h0681;
		end
		32'h0000A748: begin
				q			<=			16'h0097;
		end
		32'h0000A74A: begin
				q			<=			16'h0000;
		end
		32'h0000A74C: begin
				q			<=			16'h80E7;
		end
		32'h0000A74E: begin
				q			<=			16'hE280;
		end
		32'h0000A750: begin
				q			<=			16'h0413;
		end
		32'h0000A752: begin
				q			<=			16'h0005;
		end
		32'h0000A754: begin
				q			<=			16'h0593;
		end
		32'h0000A756: begin
				q			<=			16'h0081;
		end
		32'h0000A758: begin
				q			<=			16'h8513;
		end
		32'h0000A75A: begin
				q			<=			16'h0004;
		end
		32'h0000A75C: begin
				q			<=			16'h0097;
		end
		32'h0000A75E: begin
				q			<=			16'h0000;
		end
		32'h0000A760: begin
				q			<=			16'h80E7;
		end
		32'h0000A762: begin
				q			<=			16'hD740;
		end
		32'h0000A764: begin
				q			<=			16'h0513;
		end
		32'h0000A766: begin
				q			<=			16'h0004;
		end
		32'h0000A768: begin
				q			<=			16'h2083;
		end
		32'h0000A76A: begin
				q			<=			16'h07C1;
		end
		32'h0000A76C: begin
				q			<=			16'h2403;
		end
		32'h0000A76E: begin
				q			<=			16'h0781;
		end
		32'h0000A770: begin
				q			<=			16'h2483;
		end
		32'h0000A772: begin
				q			<=			16'h0741;
		end
		32'h0000A774: begin
				q			<=			16'h0113;
		end
		32'h0000A776: begin
				q			<=			16'h0801;
		end
		32'h0000A778: begin
				q			<=			16'h8067;
		end
		32'h0000A77A: begin
				q			<=			16'h0000;
		end
		32'h0000A77C: begin
				q			<=			16'h8613;
		end
		32'h0000A77E: begin
				q			<=			16'h0005;
		end
		32'h0000A780: begin
				q			<=			16'h0713;
		end
		32'h0000A782: begin
				q			<=			16'h0000;
		end
		32'h0000A784: begin
				q			<=			16'h0593;
		end
		32'h0000A786: begin
				q			<=			16'h0005;
		end
		32'h0000A788: begin
				q			<=			16'h0693;
		end
		32'h0000A78A: begin
				q			<=			16'h0000;
		end
		32'h0000A78C: begin
				q			<=			16'h0513;
		end
		32'h0000A78E: begin
				q			<=			16'h4090;
		end
		32'h0000A790: begin
				q			<=			16'hF06F;
		end
		32'h0000A792: begin
				q			<=			16'hDE1F;
		end
		32'h0000A794: begin
				q			<=			16'h8713;
		end
		32'h0000A796: begin
				q			<=			16'h0006;
		end
		32'h0000A798: begin
				q			<=			16'h0693;
		end
		32'h0000A79A: begin
				q			<=			16'h0006;
		end
		32'h0000A79C: begin
				q			<=			16'h8613;
		end
		32'h0000A79E: begin
				q			<=			16'h0005;
		end
		32'h0000A7A0: begin
				q			<=			16'h0593;
		end
		32'h0000A7A2: begin
				q			<=			16'h0005;
		end
		32'h0000A7A4: begin
				q			<=			16'h0513;
		end
		32'h0000A7A6: begin
				q			<=			16'h0300;
		end
		32'h0000A7A8: begin
				q			<=			16'h0317;
		end
		32'h0000A7AA: begin
				q			<=			16'h0000;
		end
		32'h0000A7AC: begin
				q			<=			16'h0067;
		end
		32'h0000A7AE: begin
				q			<=			16'hDC83;
		end
		32'h0000A7B0: begin
				q			<=			16'h0593;
		end
		32'h0000A7B2: begin
				q			<=			16'h0005;
		end
		32'h0000A7B4: begin
				q			<=			16'h0713;
		end
		32'h0000A7B6: begin
				q			<=			16'h0000;
		end
		32'h0000A7B8: begin
				q			<=			16'h0693;
		end
		32'h0000A7BA: begin
				q			<=			16'h0000;
		end
		32'h0000A7BC: begin
				q			<=			16'h0613;
		end
		32'h0000A7BE: begin
				q			<=			16'h0000;
		end
		32'h0000A7C0: begin
				q			<=			16'h0513;
		end
		32'h0000A7C2: begin
				q			<=			16'h0390;
		end
		32'h0000A7C4: begin
				q			<=			16'hF06F;
		end
		32'h0000A7C6: begin
				q			<=			16'hDADF;
		end
		32'h0000A7C8: begin
				q			<=			16'h8613;
		end
		32'h0000A7CA: begin
				q			<=			16'h0005;
		end
		32'h0000A7CC: begin
				q			<=			16'h0713;
		end
		32'h0000A7CE: begin
				q			<=			16'h0000;
		end
		32'h0000A7D0: begin
				q			<=			16'h0593;
		end
		32'h0000A7D2: begin
				q			<=			16'h0005;
		end
		32'h0000A7D4: begin
				q			<=			16'h0693;
		end
		32'h0000A7D6: begin
				q			<=			16'h0000;
		end
		32'h0000A7D8: begin
				q			<=			16'h0513;
		end
		32'h0000A7DA: begin
				q			<=			16'h4010;
		end
		32'h0000A7DC: begin
				q			<=			16'h0317;
		end
		32'h0000A7DE: begin
				q			<=			16'h0000;
		end
		32'h0000A7E0: begin
				q			<=			16'h0067;
		end
		32'h0000A7E2: begin
				q			<=			16'hD943;
		end
		32'h0000A7E4: begin
				q			<=			16'h0593;
		end
		32'h0000A7E6: begin
				q			<=			16'h0005;
		end
		32'h0000A7E8: begin
				q			<=			16'h0713;
		end
		32'h0000A7EA: begin
				q			<=			16'h0000;
		end
		32'h0000A7EC: begin
				q			<=			16'h0693;
		end
		32'h0000A7EE: begin
				q			<=			16'h0000;
		end
		32'h0000A7F0: begin
				q			<=			16'h0613;
		end
		32'h0000A7F2: begin
				q			<=			16'h0000;
		end
		32'h0000A7F4: begin
				q			<=			16'h0513;
		end
		32'h0000A7F6: begin
				q			<=			16'h4020;
		end
		32'h0000A7F8: begin
				q			<=			16'hF06F;
		end
		32'h0000A7FA: begin
				q			<=			16'hD79F;
		end
		32'h0000A7FC: begin
				q			<=			16'h0113;
		end
		32'h0000A7FE: begin
				q			<=			16'hFF01;
		end
		32'h0000A800: begin
				q			<=			16'h2623;
		end
		32'h0000A802: begin
				q			<=			16'h0011;
		end
		32'h0000A804: begin
				q			<=			16'h0097;
		end
		32'h0000A806: begin
				q			<=			16'h0000;
		end
		32'h0000A808: begin
				q			<=			16'h80E7;
		end
		32'h0000A80A: begin
				q			<=			16'h2940;
		end
		32'h0000A80C: begin
				q			<=			16'h2083;
		end
		32'h0000A80E: begin
				q			<=			16'h00C1;
		end
		32'h0000A810: begin
				q			<=			16'h0793;
		end
		32'h0000A812: begin
				q			<=			16'h00C0;
		end
		32'h0000A814: begin
				q			<=			16'h2023;
		end
		32'h0000A816: begin
				q			<=			16'h00F5;
		end
		32'h0000A818: begin
				q			<=			16'h0513;
		end
		32'h0000A81A: begin
				q			<=			16'hFFF0;
		end
		32'h0000A81C: begin
				q			<=			16'h0113;
		end
		32'h0000A81E: begin
				q			<=			16'h0101;
		end
		32'h0000A820: begin
				q			<=			16'h8067;
		end
		32'h0000A822: begin
				q			<=			16'h0000;
		end
		32'h0000A824: begin
				q			<=			16'h0113;
		end
		32'h0000A826: begin
				q			<=			16'hFF01;
		end
		32'h0000A828: begin
				q			<=			16'h2623;
		end
		32'h0000A82A: begin
				q			<=			16'h0011;
		end
		32'h0000A82C: begin
				q			<=			16'h00EF;
		end
		32'h0000A82E: begin
				q			<=			16'h26C0;
		end
		32'h0000A830: begin
				q			<=			16'h2083;
		end
		32'h0000A832: begin
				q			<=			16'h00C1;
		end
		32'h0000A834: begin
				q			<=			16'h0793;
		end
		32'h0000A836: begin
				q			<=			16'h00B0;
		end
		32'h0000A838: begin
				q			<=			16'h2023;
		end
		32'h0000A83A: begin
				q			<=			16'h00F5;
		end
		32'h0000A83C: begin
				q			<=			16'h0513;
		end
		32'h0000A83E: begin
				q			<=			16'hFFF0;
		end
		32'h0000A840: begin
				q			<=			16'h0113;
		end
		32'h0000A842: begin
				q			<=			16'h0101;
		end
		32'h0000A844: begin
				q			<=			16'h8067;
		end
		32'h0000A846: begin
				q			<=			16'h0000;
		end
		32'h0000A848: begin
				q			<=			16'h0513;
		end
		32'h0000A84A: begin
				q			<=			16'h0010;
		end
		32'h0000A84C: begin
				q			<=			16'h8067;
		end
		32'h0000A84E: begin
				q			<=			16'h0000;
		end
		32'h0000A850: begin
				q			<=			16'h0113;
		end
		32'h0000A852: begin
				q			<=			16'hFF01;
		end
		32'h0000A854: begin
				q			<=			16'h2623;
		end
		32'h0000A856: begin
				q			<=			16'h0011;
		end
		32'h0000A858: begin
				q			<=			16'h00EF;
		end
		32'h0000A85A: begin
				q			<=			16'h2400;
		end
		32'h0000A85C: begin
				q			<=			16'h2083;
		end
		32'h0000A85E: begin
				q			<=			16'h00C1;
		end
		32'h0000A860: begin
				q			<=			16'h0793;
		end
		32'h0000A862: begin
				q			<=			16'h0160;
		end
		32'h0000A864: begin
				q			<=			16'h2023;
		end
		32'h0000A866: begin
				q			<=			16'h00F5;
		end
		32'h0000A868: begin
				q			<=			16'h0513;
		end
		32'h0000A86A: begin
				q			<=			16'hFFF0;
		end
		32'h0000A86C: begin
				q			<=			16'h0113;
		end
		32'h0000A86E: begin
				q			<=			16'h0101;
		end
		32'h0000A870: begin
				q			<=			16'h8067;
		end
		32'h0000A872: begin
				q			<=			16'h0000;
		end
		32'h0000A874: begin
				q			<=			16'h0113;
		end
		32'h0000A876: begin
				q			<=			16'hFF01;
		end
		32'h0000A878: begin
				q			<=			16'h2623;
		end
		32'h0000A87A: begin
				q			<=			16'h0011;
		end
		32'h0000A87C: begin
				q			<=			16'h0097;
		end
		32'h0000A87E: begin
				q			<=			16'h0000;
		end
		32'h0000A880: begin
				q			<=			16'h80E7;
		end
		32'h0000A882: begin
				q			<=			16'h21C0;
		end
		32'h0000A884: begin
				q			<=			16'h2083;
		end
		32'h0000A886: begin
				q			<=			16'h00C1;
		end
		32'h0000A888: begin
				q			<=			16'h0793;
		end
		32'h0000A88A: begin
				q			<=			16'h00A0;
		end
		32'h0000A88C: begin
				q			<=			16'h2023;
		end
		32'h0000A88E: begin
				q			<=			16'h00F5;
		end
		32'h0000A890: begin
				q			<=			16'h0513;
		end
		32'h0000A892: begin
				q			<=			16'hFFF0;
		end
		32'h0000A894: begin
				q			<=			16'h0113;
		end
		32'h0000A896: begin
				q			<=			16'h0101;
		end
		32'h0000A898: begin
				q			<=			16'h8067;
		end
		32'h0000A89A: begin
				q			<=			16'h0000;
		end
		32'h0000A89C: begin
				q			<=			16'h0113;
		end
		32'h0000A89E: begin
				q			<=			16'hFB01;
		end
		32'h0000A8A0: begin
				q			<=			16'h0593;
		end
		32'h0000A8A2: begin
				q			<=			16'h0041;
		end
		32'h0000A8A4: begin
				q			<=			16'h2623;
		end
		32'h0000A8A6: begin
				q			<=			16'h0411;
		end
		32'h0000A8A8: begin
				q			<=			16'hF0EF;
		end
		32'h0000A8AA: begin
				q			<=			16'hD75F;
		end
		32'h0000A8AC: begin
				q			<=			16'h0793;
		end
		32'h0000A8AE: begin
				q			<=			16'hFFF0;
		end
		32'h0000A8B0: begin
				q			<=			16'h0863;
		end
		32'h0000A8B2: begin
				q			<=			16'h00F5;
		end
		32'h0000A8B4: begin
				q			<=			16'h2503;
		end
		32'h0000A8B6: begin
				q			<=			16'h0081;
		end
		32'h0000A8B8: begin
				q			<=			16'h5513;
		end
		32'h0000A8BA: begin
				q			<=			16'h00D5;
		end
		32'h0000A8BC: begin
				q			<=			16'h7513;
		end
		32'h0000A8BE: begin
				q			<=			16'h0015;
		end
		32'h0000A8C0: begin
				q			<=			16'h2083;
		end
		32'h0000A8C2: begin
				q			<=			16'h04C1;
		end
		32'h0000A8C4: begin
				q			<=			16'h0113;
		end
		32'h0000A8C6: begin
				q			<=			16'h0501;
		end
		32'h0000A8C8: begin
				q			<=			16'h8067;
		end
		32'h0000A8CA: begin
				q			<=			16'h0000;
		end
		32'h0000A8CC: begin
				q			<=			16'h0593;
		end
		32'h0000A8CE: begin
				q			<=			16'h0005;
		end
		32'h0000A8D0: begin
				q			<=			16'h0713;
		end
		32'h0000A8D2: begin
				q			<=			16'h0000;
		end
		32'h0000A8D4: begin
				q			<=			16'h0693;
		end
		32'h0000A8D6: begin
				q			<=			16'h0000;
		end
		32'h0000A8D8: begin
				q			<=			16'h0613;
		end
		32'h0000A8DA: begin
				q			<=			16'h0000;
		end
		32'h0000A8DC: begin
				q			<=			16'h0513;
		end
		32'h0000A8DE: begin
				q			<=			16'h0A90;
		end
		32'h0000A8E0: begin
				q			<=			16'h0317;
		end
		32'h0000A8E2: begin
				q			<=			16'h0000;
		end
		32'h0000A8E4: begin
				q			<=			16'h0067;
		end
		32'h0000A8E6: begin
				q			<=			16'hC903;
		end
		32'h0000A8E8: begin
				q			<=			16'h0113;
		end
		32'h0000A8EA: begin
				q			<=			16'hFE01;
		end
		32'h0000A8EC: begin
				q			<=			16'h2C23;
		end
		32'h0000A8EE: begin
				q			<=			16'h0081;
		end
		32'h0000A8F0: begin
				q			<=			16'h6417;
		end
		32'h0000A8F2: begin
				q			<=			16'h0000;
		end
		32'h0000A8F4: begin
				q			<=			16'h0413;
		end
		32'h0000A8F6: begin
				q			<=			16'h6C44;
		end
		32'h0000A8F8: begin
				q			<=			16'h2783;
		end
		32'h0000A8FA: begin
				q			<=			16'h0004;
		end
		32'h0000A8FC: begin
				q			<=			16'h2A23;
		end
		32'h0000A8FE: begin
				q			<=			16'h0091;
		end
		32'h0000A900: begin
				q			<=			16'h2E23;
		end
		32'h0000A902: begin
				q			<=			16'h0011;
		end
		32'h0000A904: begin
				q			<=			16'h0493;
		end
		32'h0000A906: begin
				q			<=			16'h0005;
		end
		32'h0000A908: begin
				q			<=			16'h9A63;
		end
		32'h0000A90A: begin
				q			<=			16'h0007;
		end
		32'h0000A90C: begin
				q			<=			16'h0593;
		end
		32'h0000A90E: begin
				q			<=			16'h0000;
		end
		32'h0000A910: begin
				q			<=			16'h0513;
		end
		32'h0000A912: begin
				q			<=			16'h0004;
		end
		32'h0000A914: begin
				q			<=			16'h0097;
		end
		32'h0000A916: begin
				q			<=			16'h0000;
		end
		32'h0000A918: begin
				q			<=			16'h80E7;
		end
		32'h0000A91A: begin
				q			<=			16'hFB80;
		end
		32'h0000A91C: begin
				q			<=			16'h0513;
		end
		32'h0000A91E: begin
				q			<=			16'h0081;
		end
		32'h0000A920: begin
				q			<=			16'h0593;
		end
		32'h0000A922: begin
				q			<=			16'h0000;
		end
		32'h0000A924: begin
				q			<=			16'h0097;
		end
		32'h0000A926: begin
				q			<=			16'h0000;
		end
		32'h0000A928: begin
				q			<=			16'h80E7;
		end
		32'h0000A92A: begin
				q			<=			16'hFA80;
		end
		32'h0000A92C: begin
				q			<=			16'h2703;
		end
		32'h0000A92E: begin
				q			<=			16'h0004;
		end
		32'h0000A930: begin
				q			<=			16'h2783;
		end
		32'h0000A932: begin
				q			<=			16'h0081;
		end
		32'h0000A934: begin
				q			<=			16'h2683;
		end
		32'h0000A936: begin
				q			<=			16'h0044;
		end
		32'h0000A938: begin
				q			<=			16'h2083;
		end
		32'h0000A93A: begin
				q			<=			16'h01C1;
		end
		32'h0000A93C: begin
				q			<=			16'h87B3;
		end
		32'h0000A93E: begin
				q			<=			16'h40E7;
		end
		32'h0000A940: begin
				q			<=			16'h4737;
		end
		32'h0000A942: begin
				q			<=			16'h000F;
		end
		32'h0000A944: begin
				q			<=			16'h0713;
		end
		32'h0000A946: begin
				q			<=			16'h2407;
		end
		32'h0000A948: begin
				q			<=			16'h87B3;
		end
		32'h0000A94A: begin
				q			<=			16'h02E7;
		end
		32'h0000A94C: begin
				q			<=			16'h2703;
		end
		32'h0000A94E: begin
				q			<=			16'h00C1;
		end
		32'h0000A950: begin
				q			<=			16'h2403;
		end
		32'h0000A952: begin
				q			<=			16'h0181;
		end
		32'h0000A954: begin
				q			<=			16'hA423;
		end
		32'h0000A956: begin
				q			<=			16'h0004;
		end
		32'h0000A958: begin
				q			<=			16'h0733;
		end
		32'h0000A95A: begin
				q			<=			16'h40D7;
		end
		32'h0000A95C: begin
				q			<=			16'hA623;
		end
		32'h0000A95E: begin
				q			<=			16'h0004;
		end
		32'h0000A960: begin
				q			<=			16'hA223;
		end
		32'h0000A962: begin
				q			<=			16'h0004;
		end
		32'h0000A964: begin
				q			<=			16'h0513;
		end
		32'h0000A966: begin
				q			<=			16'hFFF0;
		end
		32'h0000A968: begin
				q			<=			16'h87B3;
		end
		32'h0000A96A: begin
				q			<=			16'h00E7;
		end
		32'h0000A96C: begin
				q			<=			16'hA023;
		end
		32'h0000A96E: begin
				q			<=			16'h00F4;
		end
		32'h0000A970: begin
				q			<=			16'h2483;
		end
		32'h0000A972: begin
				q			<=			16'h0141;
		end
		32'h0000A974: begin
				q			<=			16'h0113;
		end
		32'h0000A976: begin
				q			<=			16'h0201;
		end
		32'h0000A978: begin
				q			<=			16'h8067;
		end
		32'h0000A97A: begin
				q			<=			16'h0000;
		end
		32'h0000A97C: begin
				q			<=			16'h1223;
		end
		32'h0000A97E: begin
				q			<=			16'h0005;
		end
		32'h0000A980: begin
				q			<=			16'h2023;
		end
		32'h0000A982: begin
				q			<=			16'h0005;
		end
		32'h0000A984: begin
				q			<=			16'h0513;
		end
		32'h0000A986: begin
				q			<=			16'h0000;
		end
		32'h0000A988: begin
				q			<=			16'h8067;
		end
		32'h0000A98A: begin
				q			<=			16'h0000;
		end
		32'h0000A98C: begin
				q			<=			16'h0513;
		end
		32'h0000A98E: begin
				q			<=			16'hFFF0;
		end
		32'h0000A990: begin
				q			<=			16'h8067;
		end
		32'h0000A992: begin
				q			<=			16'h0000;
		end
		32'h0000A994: begin
				q			<=			16'h0513;
		end
		32'h0000A996: begin
				q			<=			16'hFFF0;
		end
		32'h0000A998: begin
				q			<=			16'h8067;
		end
		32'h0000A99A: begin
				q			<=			16'h0000;
		end
		32'h0000A99C: begin
				q			<=			16'h0513;
		end
		32'h0000A99E: begin
				q			<=			16'hFFF0;
		end
		32'h0000A9A0: begin
				q			<=			16'h8067;
		end
		32'h0000A9A2: begin
				q			<=			16'h0000;
		end
		32'h0000A9A4: begin
				q			<=			16'h0513;
		end
		32'h0000A9A6: begin
				q			<=			16'hFFF0;
		end
		32'h0000A9A8: begin
				q			<=			16'h8067;
		end
		32'h0000A9AA: begin
				q			<=			16'h0000;
		end
		32'h0000A9AC: begin
				q			<=			16'h0513;
		end
		32'h0000A9AE: begin
				q			<=			16'h0000;
		end
		32'h0000A9B0: begin
				q			<=			16'h8067;
		end
		32'h0000A9B2: begin
				q			<=			16'h0000;
		end
		32'h0000A9B4: begin
				q			<=			16'h0793;
		end
		32'h0000A9B6: begin
				q			<=			16'h0020;
		end
		32'h0000A9B8: begin
				q			<=			16'h0663;
		end
		32'h0000A9BA: begin
				q			<=			16'h00F5;
		end
		32'h0000A9BC: begin
				q			<=			16'h0513;
		end
		32'h0000A9BE: begin
				q			<=			16'hFFF0;
		end
		32'h0000A9C0: begin
				q			<=			16'h8067;
		end
		32'h0000A9C2: begin
				q			<=			16'h0000;
		end
		32'h0000A9C4: begin
				q			<=			16'h4537;
		end
		32'h0000A9C6: begin
				q			<=			16'h000F;
		end
		32'h0000A9C8: begin
				q			<=			16'h0513;
		end
		32'h0000A9CA: begin
				q			<=			16'h2405;
		end
		32'h0000A9CC: begin
				q			<=			16'h8067;
		end
		32'h0000A9CE: begin
				q			<=			16'h0000;
		end
		32'h0000A9D0: begin
				q			<=			16'h0113;
		end
		32'h0000A9D2: begin
				q			<=			16'hFF01;
		end
		32'h0000A9D4: begin
				q			<=			16'h2423;
		end
		32'h0000A9D6: begin
				q			<=			16'h0081;
		end
		32'h0000A9D8: begin
				q			<=			16'h6417;
		end
		32'h0000A9DA: begin
				q			<=			16'h0000;
		end
		32'h0000A9DC: begin
				q			<=			16'h0413;
		end
		32'h0000A9DE: begin
				q			<=			16'h5D84;
		end
		32'h0000A9E0: begin
				q			<=			16'h2783;
		end
		32'h0000A9E2: begin
				q			<=			16'h0004;
		end
		32'h0000A9E4: begin
				q			<=			16'h2223;
		end
		32'h0000A9E6: begin
				q			<=			16'h0091;
		end
		32'h0000A9E8: begin
				q			<=			16'h2623;
		end
		32'h0000A9EA: begin
				q			<=			16'h0011;
		end
		32'h0000A9EC: begin
				q			<=			16'h0493;
		end
		32'h0000A9EE: begin
				q			<=			16'h0005;
		end
		32'h0000A9F0: begin
				q			<=			16'h9263;
		end
		32'h0000A9F2: begin
				q			<=			16'h0407;
		end
		32'h0000A9F4: begin
				q			<=			16'h0713;
		end
		32'h0000A9F6: begin
				q			<=			16'h0000;
		end
		32'h0000A9F8: begin
				q			<=			16'h0693;
		end
		32'h0000A9FA: begin
				q			<=			16'h0000;
		end
		32'h0000A9FC: begin
				q			<=			16'h0613;
		end
		32'h0000A9FE: begin
				q			<=			16'h0000;
		end
		32'h0000AA00: begin
				q			<=			16'h0593;
		end
		32'h0000AA02: begin
				q			<=			16'h0000;
		end
		32'h0000AA04: begin
				q			<=			16'h0513;
		end
		32'h0000AA06: begin
				q			<=			16'h0D60;
		end
		32'h0000AA08: begin
				q			<=			16'hF0EF;
		end
		32'h0000AA0A: begin
				q			<=			16'hB69F;
		end
		32'h0000AA0C: begin
				q			<=			16'h0793;
		end
		32'h0000AA0E: begin
				q			<=			16'hFFF0;
		end
		32'h0000AA10: begin
				q			<=			16'h1E63;
		end
		32'h0000AA12: begin
				q			<=			16'h00F5;
		end
		32'h0000AA14: begin
				q			<=			16'h0513;
		end
		32'h0000AA16: begin
				q			<=			16'hFFF0;
		end
		32'h0000AA18: begin
				q			<=			16'h2083;
		end
		32'h0000AA1A: begin
				q			<=			16'h00C1;
		end
		32'h0000AA1C: begin
				q			<=			16'h2403;
		end
		32'h0000AA1E: begin
				q			<=			16'h0081;
		end
		32'h0000AA20: begin
				q			<=			16'h2483;
		end
		32'h0000AA22: begin
				q			<=			16'h0041;
		end
		32'h0000AA24: begin
				q			<=			16'h0113;
		end
		32'h0000AA26: begin
				q			<=			16'h0101;
		end
		32'h0000AA28: begin
				q			<=			16'h8067;
		end
		32'h0000AA2A: begin
				q			<=			16'h0000;
		end
		32'h0000AA2C: begin
				q			<=			16'h6797;
		end
		32'h0000AA2E: begin
				q			<=			16'h0000;
		end
		32'h0000AA30: begin
				q			<=			16'hA223;
		end
		32'h0000AA32: begin
				q			<=			16'h58A7;
		end
		32'h0000AA34: begin
				q			<=			16'h2583;
		end
		32'h0000AA36: begin
				q			<=			16'h0004;
		end
		32'h0000AA38: begin
				q			<=			16'h0713;
		end
		32'h0000AA3A: begin
				q			<=			16'h0000;
		end
		32'h0000AA3C: begin
				q			<=			16'h0693;
		end
		32'h0000AA3E: begin
				q			<=			16'h0000;
		end
		32'h0000AA40: begin
				q			<=			16'h85B3;
		end
		32'h0000AA42: begin
				q			<=			16'h00B4;
		end
		32'h0000AA44: begin
				q			<=			16'h0613;
		end
		32'h0000AA46: begin
				q			<=			16'h0000;
		end
		32'h0000AA48: begin
				q			<=			16'h0513;
		end
		32'h0000AA4A: begin
				q			<=			16'h0D60;
		end
		32'h0000AA4C: begin
				q			<=			16'hF0EF;
		end
		32'h0000AA4E: begin
				q			<=			16'hB25F;
		end
		32'h0000AA50: begin
				q			<=			16'h2783;
		end
		32'h0000AA52: begin
				q			<=			16'h0004;
		end
		32'h0000AA54: begin
				q			<=			16'h84B3;
		end
		32'h0000AA56: begin
				q			<=			16'h00F4;
		end
		32'h0000AA58: begin
				q			<=			16'h1EE3;
		end
		32'h0000AA5A: begin
				q			<=			16'hFA95;
		end
		32'h0000AA5C: begin
				q			<=			16'h6717;
		end
		32'h0000AA5E: begin
				q			<=			16'h0000;
		end
		32'h0000AA60: begin
				q			<=			16'h2A23;
		end
		32'h0000AA62: begin
				q			<=			16'h54A7;
		end
		32'h0000AA64: begin
				q			<=			16'h8513;
		end
		32'h0000AA66: begin
				q			<=			16'h0007;
		end
		32'h0000AA68: begin
				q			<=			16'hF06F;
		end
		32'h0000AA6A: begin
				q			<=			16'hFB1F;
		end
		32'h0000AA6C: begin
				q			<=			16'h0113;
		end
		32'h0000AA6E: begin
				q			<=			16'hFF01;
		end
		32'h0000AA70: begin
				q			<=			16'h0593;
		end
		32'h0000AA72: begin
				q			<=			16'h0005;
		end
		32'h0000AA74: begin
				q			<=			16'h0713;
		end
		32'h0000AA76: begin
				q			<=			16'h0000;
		end
		32'h0000AA78: begin
				q			<=			16'h0693;
		end
		32'h0000AA7A: begin
				q			<=			16'h0000;
		end
		32'h0000AA7C: begin
				q			<=			16'h0613;
		end
		32'h0000AA7E: begin
				q			<=			16'h0000;
		end
		32'h0000AA80: begin
				q			<=			16'h0513;
		end
		32'h0000AA82: begin
				q			<=			16'h05D0;
		end
		32'h0000AA84: begin
				q			<=			16'h2623;
		end
		32'h0000AA86: begin
				q			<=			16'h0011;
		end
		32'h0000AA88: begin
				q			<=			16'h0097;
		end
		32'h0000AA8A: begin
				q			<=			16'h0000;
		end
		32'h0000AA8C: begin
				q			<=			16'h80E7;
		end
		32'h0000AA8E: begin
				q			<=			16'hAE80;
		end
		32'h0000AA90: begin
				q			<=			16'h006F;
		end
		32'h0000AA92: begin
				q			<=			16'h0000;
		end
		32'h0000AA94: begin
				q			<=			16'h0000;
		end
		32'h0000AA96: begin
				q			<=			16'h0000;
		end
		32'h0000AA98: begin
				q			<=			16'h6797;
		end
		32'h0000AA9A: begin
				q			<=			16'h0000;
		end
		32'h0000AA9C: begin
				q			<=			16'h8793;
		end
		32'h0000AA9E: begin
				q			<=			16'hE407;
		end
		32'h0000AAA0: begin
				q			<=			16'hA503;
		end
		32'h0000AAA2: begin
				q			<=			16'h0007;
		end
		32'h0000AAA4: begin
				q			<=			16'h8067;
		end
		32'h0000AAA6: begin
				q			<=			16'h0000;
		end
		32'h0000AAA8: begin
				q			<=			16'h0000;
		end
		32'h0000AAAA: begin
				q			<=			16'h0000;
		end
		32'h0000AAAC: begin
				q			<=			16'h8793;
		end
		32'h0000AAAE: begin
				q			<=			16'h0005;
		end
		32'h0000AAB0: begin
				q			<=			16'h0813;
		end
		32'h0000AAB2: begin
				q			<=			16'h0006;
		end
		32'h0000AAB4: begin
				q			<=			16'h8713;
		end
		32'h0000AAB6: begin
				q			<=			16'h0006;
		end
		32'h0000AAB8: begin
				q			<=			16'h0313;
		end
		32'h0000AABA: begin
				q			<=			16'h0005;
		end
		32'h0000AABC: begin
				q			<=			16'h9663;
		end
		32'h0000AABE: begin
				q			<=			16'h2806;
		end
		32'h0000AAC0: begin
				q			<=			16'h5897;
		end
		32'h0000AAC2: begin
				q			<=			16'h0000;
		end
		32'h0000AAC4: begin
				q			<=			16'h8893;
		end
		32'h0000AAC6: begin
				q			<=			16'hEAC8;
		end
		32'h0000AAC8: begin
				q			<=			16'hF663;
		end
		32'h0000AACA: begin
				q			<=			16'h0EC5;
		end
		32'h0000AACC: begin
				q			<=			16'h0737;
		end
		32'h0000AACE: begin
				q			<=			16'h0001;
		end
		32'h0000AAD0: begin
				q			<=			16'h7863;
		end
		32'h0000AAD2: begin
				q			<=			16'h0CE6;
		end
		32'h0000AAD4: begin
				q			<=			16'h0713;
		end
		32'h0000AAD6: begin
				q			<=			16'h0FF0;
		end
		32'h0000AAD8: begin
				q			<=			16'h3733;
		end
		32'h0000AADA: begin
				q			<=			16'h00C7;
		end
		32'h0000AADC: begin
				q			<=			16'h1713;
		end
		32'h0000AADE: begin
				q			<=			16'h0037;
		end
		32'h0000AAE0: begin
				q			<=			16'h56B3;
		end
		32'h0000AAE2: begin
				q			<=			16'h00E6;
		end
		32'h0000AAE4: begin
				q			<=			16'h88B3;
		end
		32'h0000AAE6: begin
				q			<=			16'h00D8;
		end
		32'h0000AAE8: begin
				q			<=			16'hC683;
		end
		32'h0000AAEA: begin
				q			<=			16'h0008;
		end
		32'h0000AAEC: begin
				q			<=			16'h8733;
		end
		32'h0000AAEE: begin
				q			<=			16'h00E6;
		end
		32'h0000AAF0: begin
				q			<=			16'h0693;
		end
		32'h0000AAF2: begin
				q			<=			16'h0200;
		end
		32'h0000AAF4: begin
				q			<=			16'h86B3;
		end
		32'h0000AAF6: begin
				q			<=			16'h40E6;
		end
		32'h0000AAF8: begin
				q			<=			16'h8C63;
		end
		32'h0000AAFA: begin
				q			<=			16'h0006;
		end
		32'h0000AAFC: begin
				q			<=			16'h97B3;
		end
		32'h0000AAFE: begin
				q			<=			16'h00D7;
		end
		32'h0000AB00: begin
				q			<=			16'h5733;
		end
		32'h0000AB02: begin
				q			<=			16'h00E5;
		end
		32'h0000AB04: begin
				q			<=			16'h1833;
		end
		32'h0000AB06: begin
				q			<=			16'h00D6;
		end
		32'h0000AB08: begin
				q			<=			16'h65B3;
		end
		32'h0000AB0A: begin
				q			<=			16'h00F7;
		end
		32'h0000AB0C: begin
				q			<=			16'h1333;
		end
		32'h0000AB0E: begin
				q			<=			16'h00D5;
		end
		32'h0000AB10: begin
				q			<=			16'h5513;
		end
		32'h0000AB12: begin
				q			<=			16'h0108;
		end
		32'h0000AB14: begin
				q			<=			16'hD7B3;
		end
		32'h0000AB16: begin
				q			<=			16'h02A5;
		end
		32'h0000AB18: begin
				q			<=			16'h1613;
		end
		32'h0000AB1A: begin
				q			<=			16'h0108;
		end
		32'h0000AB1C: begin
				q			<=			16'h5613;
		end
		32'h0000AB1E: begin
				q			<=			16'h0106;
		end
		32'h0000AB20: begin
				q			<=			16'h5693;
		end
		32'h0000AB22: begin
				q			<=			16'h0103;
		end
		32'h0000AB24: begin
				q			<=			16'hF733;
		end
		32'h0000AB26: begin
				q			<=			16'h02A5;
		end
		32'h0000AB28: begin
				q			<=			16'h05B3;
		end
		32'h0000AB2A: begin
				q			<=			16'h02F6;
		end
		32'h0000AB2C: begin
				q			<=			16'h1713;
		end
		32'h0000AB2E: begin
				q			<=			16'h0107;
		end
		32'h0000AB30: begin
				q			<=			16'h66B3;
		end
		32'h0000AB32: begin
				q			<=			16'h00D7;
		end
		32'h0000AB34: begin
				q			<=			16'h8713;
		end
		32'h0000AB36: begin
				q			<=			16'h0007;
		end
		32'h0000AB38: begin
				q			<=			16'hFE63;
		end
		32'h0000AB3A: begin
				q			<=			16'h00B6;
		end
		32'h0000AB3C: begin
				q			<=			16'h86B3;
		end
		32'h0000AB3E: begin
				q			<=			16'h0106;
		end
		32'h0000AB40: begin
				q			<=			16'h8713;
		end
		32'h0000AB42: begin
				q			<=			16'hFFF7;
		end
		32'h0000AB44: begin
				q			<=			16'hE863;
		end
		32'h0000AB46: begin
				q			<=			16'h0106;
		end
		32'h0000AB48: begin
				q			<=			16'hF663;
		end
		32'h0000AB4A: begin
				q			<=			16'h00B6;
		end
		32'h0000AB4C: begin
				q			<=			16'h8713;
		end
		32'h0000AB4E: begin
				q			<=			16'hFFE7;
		end
		32'h0000AB50: begin
				q			<=			16'h86B3;
		end
		32'h0000AB52: begin
				q			<=			16'h0106;
		end
		32'h0000AB54: begin
				q			<=			16'h86B3;
		end
		32'h0000AB56: begin
				q			<=			16'h40B6;
		end
		32'h0000AB58: begin
				q			<=			16'hF7B3;
		end
		32'h0000AB5A: begin
				q			<=			16'h02A6;
		end
		32'h0000AB5C: begin
				q			<=			16'h1313;
		end
		32'h0000AB5E: begin
				q			<=			16'h0103;
		end
		32'h0000AB60: begin
				q			<=			16'h5313;
		end
		32'h0000AB62: begin
				q			<=			16'h0103;
		end
		32'h0000AB64: begin
				q			<=			16'hD6B3;
		end
		32'h0000AB66: begin
				q			<=			16'h02A6;
		end
		32'h0000AB68: begin
				q			<=			16'h9793;
		end
		32'h0000AB6A: begin
				q			<=			16'h0107;
		end
		32'h0000AB6C: begin
				q			<=			16'hE333;
		end
		32'h0000AB6E: begin
				q			<=			16'h0067;
		end
		32'h0000AB70: begin
				q			<=			16'h05B3;
		end
		32'h0000AB72: begin
				q			<=			16'h02D6;
		end
		32'h0000AB74: begin
				q			<=			16'h8513;
		end
		32'h0000AB76: begin
				q			<=			16'h0006;
		end
		32'h0000AB78: begin
				q			<=			16'h7C63;
		end
		32'h0000AB7A: begin
				q			<=			16'h00B3;
		end
		32'h0000AB7C: begin
				q			<=			16'h0333;
		end
		32'h0000AB7E: begin
				q			<=			16'h0068;
		end
		32'h0000AB80: begin
				q			<=			16'h8513;
		end
		32'h0000AB82: begin
				q			<=			16'hFFF6;
		end
		32'h0000AB84: begin
				q			<=			16'h6663;
		end
		32'h0000AB86: begin
				q			<=			16'h0103;
		end
		32'h0000AB88: begin
				q			<=			16'h7463;
		end
		32'h0000AB8A: begin
				q			<=			16'h00B3;
		end
		32'h0000AB8C: begin
				q			<=			16'h8513;
		end
		32'h0000AB8E: begin
				q			<=			16'hFFE6;
		end
		32'h0000AB90: begin
				q			<=			16'h1713;
		end
		32'h0000AB92: begin
				q			<=			16'h0107;
		end
		32'h0000AB94: begin
				q			<=			16'h6733;
		end
		32'h0000AB96: begin
				q			<=			16'h00A7;
		end
		32'h0000AB98: begin
				q			<=			16'h0593;
		end
		32'h0000AB9A: begin
				q			<=			16'h0000;
		end
		32'h0000AB9C: begin
				q			<=			16'h006F;
		end
		32'h0000AB9E: begin
				q			<=			16'h0E40;
		end
		32'h0000ABA0: begin
				q			<=			16'h06B7;
		end
		32'h0000ABA2: begin
				q			<=			16'h0100;
		end
		32'h0000ABA4: begin
				q			<=			16'h0713;
		end
		32'h0000ABA6: begin
				q			<=			16'h0100;
		end
		32'h0000ABA8: begin
				q			<=			16'h6CE3;
		end
		32'h0000ABAA: begin
				q			<=			16'hF2D6;
		end
		32'h0000ABAC: begin
				q			<=			16'h0713;
		end
		32'h0000ABAE: begin
				q			<=			16'h0180;
		end
		32'h0000ABB0: begin
				q			<=			16'hF06F;
		end
		32'h0000ABB2: begin
				q			<=			16'hF31F;
		end
		32'h0000ABB4: begin
				q			<=			16'h1663;
		end
		32'h0000ABB6: begin
				q			<=			16'h0006;
		end
		32'h0000ABB8: begin
				q			<=			16'h0693;
		end
		32'h0000ABBA: begin
				q			<=			16'h0010;
		end
		32'h0000ABBC: begin
				q			<=			16'hD833;
		end
		32'h0000ABBE: begin
				q			<=			16'h02C6;
		end
		32'h0000ABC0: begin
				q			<=			16'h06B7;
		end
		32'h0000ABC2: begin
				q			<=			16'h0001;
		end
		32'h0000ABC4: begin
				q			<=			16'h7263;
		end
		32'h0000ABC6: begin
				q			<=			16'h0CD8;
		end
		32'h0000ABC8: begin
				q			<=			16'h0693;
		end
		32'h0000ABCA: begin
				q			<=			16'h0FF0;
		end
		32'h0000ABCC: begin
				q			<=			16'hF463;
		end
		32'h0000ABCE: begin
				q			<=			16'h0106;
		end
		32'h0000ABD0: begin
				q			<=			16'h0713;
		end
		32'h0000ABD2: begin
				q			<=			16'h0080;
		end
		32'h0000ABD4: begin
				q			<=			16'h56B3;
		end
		32'h0000ABD6: begin
				q			<=			16'h00E8;
		end
		32'h0000ABD8: begin
				q			<=			16'h88B3;
		end
		32'h0000ABDA: begin
				q			<=			16'h00D8;
		end
		32'h0000ABDC: begin
				q			<=			16'hC683;
		end
		32'h0000ABDE: begin
				q			<=			16'h0008;
		end
		32'h0000ABE0: begin
				q			<=			16'h86B3;
		end
		32'h0000ABE2: begin
				q			<=			16'h00E6;
		end
		32'h0000ABE4: begin
				q			<=			16'h0713;
		end
		32'h0000ABE6: begin
				q			<=			16'h0200;
		end
		32'h0000ABE8: begin
				q			<=			16'h0733;
		end
		32'h0000ABEA: begin
				q			<=			16'h40D7;
		end
		32'h0000ABEC: begin
				q			<=			16'h1863;
		end
		32'h0000ABEE: begin
				q			<=			16'h0A07;
		end
		32'h0000ABF0: begin
				q			<=			16'h87B3;
		end
		32'h0000ABF2: begin
				q			<=			16'h4107;
		end
		32'h0000ABF4: begin
				q			<=			16'h0593;
		end
		32'h0000ABF6: begin
				q			<=			16'h0010;
		end
		32'h0000ABF8: begin
				q			<=			16'h5613;
		end
		32'h0000ABFA: begin
				q			<=			16'h0108;
		end
		32'h0000ABFC: begin
				q			<=			16'h1893;
		end
		32'h0000ABFE: begin
				q			<=			16'h0108;
		end
		32'h0000AC00: begin
				q			<=			16'hD893;
		end
		32'h0000AC02: begin
				q			<=			16'h0108;
		end
		32'h0000AC04: begin
				q			<=			16'h5693;
		end
		32'h0000AC06: begin
				q			<=			16'h0103;
		end
		32'h0000AC08: begin
				q			<=			16'hF733;
		end
		32'h0000AC0A: begin
				q			<=			16'h02C7;
		end
		32'h0000AC0C: begin
				q			<=			16'hD7B3;
		end
		32'h0000AC0E: begin
				q			<=			16'h02C7;
		end
		32'h0000AC10: begin
				q			<=			16'h1713;
		end
		32'h0000AC12: begin
				q			<=			16'h0107;
		end
		32'h0000AC14: begin
				q			<=			16'h66B3;
		end
		32'h0000AC16: begin
				q			<=			16'h00D7;
		end
		32'h0000AC18: begin
				q			<=			16'h8533;
		end
		32'h0000AC1A: begin
				q			<=			16'h02F8;
		end
		32'h0000AC1C: begin
				q			<=			16'h8713;
		end
		32'h0000AC1E: begin
				q			<=			16'h0007;
		end
		32'h0000AC20: begin
				q			<=			16'hFE63;
		end
		32'h0000AC22: begin
				q			<=			16'h00A6;
		end
		32'h0000AC24: begin
				q			<=			16'h86B3;
		end
		32'h0000AC26: begin
				q			<=			16'h0106;
		end
		32'h0000AC28: begin
				q			<=			16'h8713;
		end
		32'h0000AC2A: begin
				q			<=			16'hFFF7;
		end
		32'h0000AC2C: begin
				q			<=			16'hE863;
		end
		32'h0000AC2E: begin
				q			<=			16'h0106;
		end
		32'h0000AC30: begin
				q			<=			16'hF663;
		end
		32'h0000AC32: begin
				q			<=			16'h00A6;
		end
		32'h0000AC34: begin
				q			<=			16'h8713;
		end
		32'h0000AC36: begin
				q			<=			16'hFFE7;
		end
		32'h0000AC38: begin
				q			<=			16'h86B3;
		end
		32'h0000AC3A: begin
				q			<=			16'h0106;
		end
		32'h0000AC3C: begin
				q			<=			16'h86B3;
		end
		32'h0000AC3E: begin
				q			<=			16'h40A6;
		end
		32'h0000AC40: begin
				q			<=			16'hF7B3;
		end
		32'h0000AC42: begin
				q			<=			16'h02C6;
		end
		32'h0000AC44: begin
				q			<=			16'h1313;
		end
		32'h0000AC46: begin
				q			<=			16'h0103;
		end
		32'h0000AC48: begin
				q			<=			16'h5313;
		end
		32'h0000AC4A: begin
				q			<=			16'h0103;
		end
		32'h0000AC4C: begin
				q			<=			16'hD6B3;
		end
		32'h0000AC4E: begin
				q			<=			16'h02C6;
		end
		32'h0000AC50: begin
				q			<=			16'h9793;
		end
		32'h0000AC52: begin
				q			<=			16'h0107;
		end
		32'h0000AC54: begin
				q			<=			16'hE333;
		end
		32'h0000AC56: begin
				q			<=			16'h0067;
		end
		32'h0000AC58: begin
				q			<=			16'h88B3;
		end
		32'h0000AC5A: begin
				q			<=			16'h02D8;
		end
		32'h0000AC5C: begin
				q			<=			16'h8513;
		end
		32'h0000AC5E: begin
				q			<=			16'h0006;
		end
		32'h0000AC60: begin
				q			<=			16'h7C63;
		end
		32'h0000AC62: begin
				q			<=			16'h0113;
		end
		32'h0000AC64: begin
				q			<=			16'h0333;
		end
		32'h0000AC66: begin
				q			<=			16'h0068;
		end
		32'h0000AC68: begin
				q			<=			16'h8513;
		end
		32'h0000AC6A: begin
				q			<=			16'hFFF6;
		end
		32'h0000AC6C: begin
				q			<=			16'h6663;
		end
		32'h0000AC6E: begin
				q			<=			16'h0103;
		end
		32'h0000AC70: begin
				q			<=			16'h7463;
		end
		32'h0000AC72: begin
				q			<=			16'h0113;
		end
		32'h0000AC74: begin
				q			<=			16'h8513;
		end
		32'h0000AC76: begin
				q			<=			16'hFFE6;
		end
		32'h0000AC78: begin
				q			<=			16'h1713;
		end
		32'h0000AC7A: begin
				q			<=			16'h0107;
		end
		32'h0000AC7C: begin
				q			<=			16'h6733;
		end
		32'h0000AC7E: begin
				q			<=			16'h00A7;
		end
		32'h0000AC80: begin
				q			<=			16'h0513;
		end
		32'h0000AC82: begin
				q			<=			16'h0007;
		end
		32'h0000AC84: begin
				q			<=			16'h8067;
		end
		32'h0000AC86: begin
				q			<=			16'h0000;
		end
		32'h0000AC88: begin
				q			<=			16'h06B7;
		end
		32'h0000AC8A: begin
				q			<=			16'h0100;
		end
		32'h0000AC8C: begin
				q			<=			16'h0713;
		end
		32'h0000AC8E: begin
				q			<=			16'h0100;
		end
		32'h0000AC90: begin
				q			<=			16'h62E3;
		end
		32'h0000AC92: begin
				q			<=			16'hF4D8;
		end
		32'h0000AC94: begin
				q			<=			16'h0713;
		end
		32'h0000AC96: begin
				q			<=			16'h0180;
		end
		32'h0000AC98: begin
				q			<=			16'hF06F;
		end
		32'h0000AC9A: begin
				q			<=			16'hF3DF;
		end
		32'h0000AC9C: begin
				q			<=			16'h1833;
		end
		32'h0000AC9E: begin
				q			<=			16'h00E8;
		end
		32'h0000ACA0: begin
				q			<=			16'hD5B3;
		end
		32'h0000ACA2: begin
				q			<=			16'h00D7;
		end
		32'h0000ACA4: begin
				q			<=			16'h1333;
		end
		32'h0000ACA6: begin
				q			<=			16'h00E5;
		end
		32'h0000ACA8: begin
				q			<=			16'h56B3;
		end
		32'h0000ACAA: begin
				q			<=			16'h00D5;
		end
		32'h0000ACAC: begin
				q			<=			16'h5513;
		end
		32'h0000ACAE: begin
				q			<=			16'h0108;
		end
		32'h0000ACB0: begin
				q			<=			16'h97B3;
		end
		32'h0000ACB2: begin
				q			<=			16'h00E7;
		end
		32'h0000ACB4: begin
				q			<=			16'hF733;
		end
		32'h0000ACB6: begin
				q			<=			16'h02A5;
		end
		32'h0000ACB8: begin
				q			<=			16'hE8B3;
		end
		32'h0000ACBA: begin
				q			<=			16'h00F6;
		end
		32'h0000ACBC: begin
				q			<=			16'h1793;
		end
		32'h0000ACBE: begin
				q			<=			16'h0108;
		end
		32'h0000ACC0: begin
				q			<=			16'hD793;
		end
		32'h0000ACC2: begin
				q			<=			16'h0107;
		end
		32'h0000ACC4: begin
				q			<=			16'hD613;
		end
		32'h0000ACC6: begin
				q			<=			16'h0108;
		end
		32'h0000ACC8: begin
				q			<=			16'hD5B3;
		end
		32'h0000ACCA: begin
				q			<=			16'h02A5;
		end
		32'h0000ACCC: begin
				q			<=			16'h1713;
		end
		32'h0000ACCE: begin
				q			<=			16'h0107;
		end
		32'h0000ACD0: begin
				q			<=			16'h6733;
		end
		32'h0000ACD2: begin
				q			<=			16'h00C7;
		end
		32'h0000ACD4: begin
				q			<=			16'h86B3;
		end
		32'h0000ACD6: begin
				q			<=			16'h02B7;
		end
		32'h0000ACD8: begin
				q			<=			16'h8613;
		end
		32'h0000ACDA: begin
				q			<=			16'h0005;
		end
		32'h0000ACDC: begin
				q			<=			16'h7E63;
		end
		32'h0000ACDE: begin
				q			<=			16'h00D7;
		end
		32'h0000ACE0: begin
				q			<=			16'h0733;
		end
		32'h0000ACE2: begin
				q			<=			16'h0107;
		end
		32'h0000ACE4: begin
				q			<=			16'h8613;
		end
		32'h0000ACE6: begin
				q			<=			16'hFFF5;
		end
		32'h0000ACE8: begin
				q			<=			16'h6863;
		end
		32'h0000ACEA: begin
				q			<=			16'h0107;
		end
		32'h0000ACEC: begin
				q			<=			16'h7663;
		end
		32'h0000ACEE: begin
				q			<=			16'h00D7;
		end
		32'h0000ACF0: begin
				q			<=			16'h8613;
		end
		32'h0000ACF2: begin
				q			<=			16'hFFE5;
		end
		32'h0000ACF4: begin
				q			<=			16'h0733;
		end
		32'h0000ACF6: begin
				q			<=			16'h0107;
		end
		32'h0000ACF8: begin
				q			<=			16'h06B3;
		end
		32'h0000ACFA: begin
				q			<=			16'h40D7;
		end
		32'h0000ACFC: begin
				q			<=			16'hF733;
		end
		32'h0000ACFE: begin
				q			<=			16'h02A6;
		end
		32'h0000AD00: begin
				q			<=			16'h9893;
		end
		32'h0000AD02: begin
				q			<=			16'h0108;
		end
		32'h0000AD04: begin
				q			<=			16'hD893;
		end
		32'h0000AD06: begin
				q			<=			16'h0108;
		end
		32'h0000AD08: begin
				q			<=			16'hD6B3;
		end
		32'h0000AD0A: begin
				q			<=			16'h02A6;
		end
		32'h0000AD0C: begin
				q			<=			16'h1713;
		end
		32'h0000AD0E: begin
				q			<=			16'h0107;
		end
		32'h0000AD10: begin
				q			<=			16'h85B3;
		end
		32'h0000AD12: begin
				q			<=			16'h02D7;
		end
		32'h0000AD14: begin
				q			<=			16'h67B3;
		end
		32'h0000AD16: begin
				q			<=			16'h0117;
		end
		32'h0000AD18: begin
				q			<=			16'h8713;
		end
		32'h0000AD1A: begin
				q			<=			16'h0006;
		end
		32'h0000AD1C: begin
				q			<=			16'hFE63;
		end
		32'h0000AD1E: begin
				q			<=			16'h00B7;
		end
		32'h0000AD20: begin
				q			<=			16'h87B3;
		end
		32'h0000AD22: begin
				q			<=			16'h0107;
		end
		32'h0000AD24: begin
				q			<=			16'h8713;
		end
		32'h0000AD26: begin
				q			<=			16'hFFF6;
		end
		32'h0000AD28: begin
				q			<=			16'hE863;
		end
		32'h0000AD2A: begin
				q			<=			16'h0107;
		end
		32'h0000AD2C: begin
				q			<=			16'hF663;
		end
		32'h0000AD2E: begin
				q			<=			16'h00B7;
		end
		32'h0000AD30: begin
				q			<=			16'h8713;
		end
		32'h0000AD32: begin
				q			<=			16'hFFE6;
		end
		32'h0000AD34: begin
				q			<=			16'h87B3;
		end
		32'h0000AD36: begin
				q			<=			16'h0107;
		end
		32'h0000AD38: begin
				q			<=			16'h87B3;
		end
		32'h0000AD3A: begin
				q			<=			16'h40B7;
		end
		32'h0000AD3C: begin
				q			<=			16'h1593;
		end
		32'h0000AD3E: begin
				q			<=			16'h0106;
		end
		32'h0000AD40: begin
				q			<=			16'hE5B3;
		end
		32'h0000AD42: begin
				q			<=			16'h00E5;
		end
		32'h0000AD44: begin
				q			<=			16'hF06F;
		end
		32'h0000AD46: begin
				q			<=			16'hEB5F;
		end
		32'h0000AD48: begin
				q			<=			16'hE663;
		end
		32'h0000AD4A: begin
				q			<=			16'h18D5;
		end
		32'h0000AD4C: begin
				q			<=			16'h0737;
		end
		32'h0000AD4E: begin
				q			<=			16'h0001;
		end
		32'h0000AD50: begin
				q			<=			16'hF463;
		end
		32'h0000AD52: begin
				q			<=			16'h04E6;
		end
		32'h0000AD54: begin
				q			<=			16'h0813;
		end
		32'h0000AD56: begin
				q			<=			16'h0FF0;
		end
		32'h0000AD58: begin
				q			<=			16'h3733;
		end
		32'h0000AD5A: begin
				q			<=			16'h00D8;
		end
		32'h0000AD5C: begin
				q			<=			16'h1713;
		end
		32'h0000AD5E: begin
				q			<=			16'h0037;
		end
		32'h0000AD60: begin
				q			<=			16'hD833;
		end
		32'h0000AD62: begin
				q			<=			16'h00E6;
		end
		32'h0000AD64: begin
				q			<=			16'h5597;
		end
		32'h0000AD66: begin
				q			<=			16'h0000;
		end
		32'h0000AD68: begin
				q			<=			16'h8593;
		end
		32'h0000AD6A: begin
				q			<=			16'hC085;
		end
		32'h0000AD6C: begin
				q			<=			16'h85B3;
		end
		32'h0000AD6E: begin
				q			<=			16'h0105;
		end
		32'h0000AD70: begin
				q			<=			16'hC803;
		end
		32'h0000AD72: begin
				q			<=			16'h0005;
		end
		32'h0000AD74: begin
				q			<=			16'h0593;
		end
		32'h0000AD76: begin
				q			<=			16'h0200;
		end
		32'h0000AD78: begin
				q			<=			16'h0833;
		end
		32'h0000AD7A: begin
				q			<=			16'h00E8;
		end
		32'h0000AD7C: begin
				q			<=			16'h85B3;
		end
		32'h0000AD7E: begin
				q			<=			16'h4105;
		end
		32'h0000AD80: begin
				q			<=			16'h9663;
		end
		32'h0000AD82: begin
				q			<=			16'h0205;
		end
		32'h0000AD84: begin
				q			<=			16'h0713;
		end
		32'h0000AD86: begin
				q			<=			16'h0010;
		end
		32'h0000AD88: begin
				q			<=			16'hECE3;
		end
		32'h0000AD8A: begin
				q			<=			16'hEEF6;
		end
		32'h0000AD8C: begin
				q			<=			16'h3533;
		end
		32'h0000AD8E: begin
				q			<=			16'h00C5;
		end
		32'h0000AD90: begin
				q			<=			16'h4713;
		end
		32'h0000AD92: begin
				q			<=			16'h0015;
		end
		32'h0000AD94: begin
				q			<=			16'hF06F;
		end
		32'h0000AD96: begin
				q			<=			16'hEEDF;
		end
		32'h0000AD98: begin
				q			<=			16'h05B7;
		end
		32'h0000AD9A: begin
				q			<=			16'h0100;
		end
		32'h0000AD9C: begin
				q			<=			16'h0713;
		end
		32'h0000AD9E: begin
				q			<=			16'h0100;
		end
		32'h0000ADA0: begin
				q			<=			16'hE0E3;
		end
		32'h0000ADA2: begin
				q			<=			16'hFCB6;
		end
		32'h0000ADA4: begin
				q			<=			16'h0713;
		end
		32'h0000ADA6: begin
				q			<=			16'h0180;
		end
		32'h0000ADA8: begin
				q			<=			16'hF06F;
		end
		32'h0000ADAA: begin
				q			<=			16'hFB9F;
		end
		32'h0000ADAC: begin
				q			<=			16'h5733;
		end
		32'h0000ADAE: begin
				q			<=			16'h0106;
		end
		32'h0000ADB0: begin
				q			<=			16'h96B3;
		end
		32'h0000ADB2: begin
				q			<=			16'h00B6;
		end
		32'h0000ADB4: begin
				q			<=			16'h66B3;
		end
		32'h0000ADB6: begin
				q			<=			16'h00D7;
		end
		32'h0000ADB8: begin
				q			<=			16'hDE93;
		end
		32'h0000ADBA: begin
				q			<=			16'h0106;
		end
		32'h0000ADBC: begin
				q			<=			16'hD733;
		end
		32'h0000ADBE: begin
				q			<=			16'h0107;
		end
		32'h0000ADC0: begin
				q			<=			16'h78B3;
		end
		32'h0000ADC2: begin
				q			<=			16'h03D7;
		end
		32'h0000ADC4: begin
				q			<=			16'h97B3;
		end
		32'h0000ADC6: begin
				q			<=			16'h00B7;
		end
		32'h0000ADC8: begin
				q			<=			16'h5833;
		end
		32'h0000ADCA: begin
				q			<=			16'h0105;
		end
		32'h0000ADCC: begin
				q			<=			16'h6333;
		end
		32'h0000ADCE: begin
				q			<=			16'h00F8;
		end
		32'h0000ADD0: begin
				q			<=			16'h9793;
		end
		32'h0000ADD2: begin
				q			<=			16'h0106;
		end
		32'h0000ADD4: begin
				q			<=			16'hD793;
		end
		32'h0000ADD6: begin
				q			<=			16'h0107;
		end
		32'h0000ADD8: begin
				q			<=			16'h5813;
		end
		32'h0000ADDA: begin
				q			<=			16'h0103;
		end
		32'h0000ADDC: begin
				q			<=			16'h1633;
		end
		32'h0000ADDE: begin
				q			<=			16'h00B6;
		end
		32'h0000ADE0: begin
				q			<=			16'h5733;
		end
		32'h0000ADE2: begin
				q			<=			16'h03D7;
		end
		32'h0000ADE4: begin
				q			<=			16'h9893;
		end
		32'h0000ADE6: begin
				q			<=			16'h0108;
		end
		32'h0000ADE8: begin
				q			<=			16'hE833;
		end
		32'h0000ADEA: begin
				q			<=			16'h0108;
		end
		32'h0000ADEC: begin
				q			<=			16'h8F33;
		end
		32'h0000ADEE: begin
				q			<=			16'h02E7;
		end
		32'h0000ADF0: begin
				q			<=			16'h0E13;
		end
		32'h0000ADF2: begin
				q			<=			16'h0007;
		end
		32'h0000ADF4: begin
				q			<=			16'h7E63;
		end
		32'h0000ADF6: begin
				q			<=			16'h01E8;
		end
		32'h0000ADF8: begin
				q			<=			16'h0833;
		end
		32'h0000ADFA: begin
				q			<=			16'h00D8;
		end
		32'h0000ADFC: begin
				q			<=			16'h0E13;
		end
		32'h0000ADFE: begin
				q			<=			16'hFFF7;
		end
		32'h0000AE00: begin
				q			<=			16'h6863;
		end
		32'h0000AE02: begin
				q			<=			16'h00D8;
		end
		32'h0000AE04: begin
				q			<=			16'h7663;
		end
		32'h0000AE06: begin
				q			<=			16'h01E8;
		end
		32'h0000AE08: begin
				q			<=			16'h0E13;
		end
		32'h0000AE0A: begin
				q			<=			16'hFFE7;
		end
		32'h0000AE0C: begin
				q			<=			16'h0833;
		end
		32'h0000AE0E: begin
				q			<=			16'h00D8;
		end
		32'h0000AE10: begin
				q			<=			16'h0833;
		end
		32'h0000AE12: begin
				q			<=			16'h41E8;
		end
		32'h0000AE14: begin
				q			<=			16'h78B3;
		end
		32'h0000AE16: begin
				q			<=			16'h03D8;
		end
		32'h0000AE18: begin
				q			<=			16'h5833;
		end
		32'h0000AE1A: begin
				q			<=			16'h03D8;
		end
		32'h0000AE1C: begin
				q			<=			16'h9893;
		end
		32'h0000AE1E: begin
				q			<=			16'h0108;
		end
		32'h0000AE20: begin
				q			<=			16'h8EB3;
		end
		32'h0000AE22: begin
				q			<=			16'h0307;
		end
		32'h0000AE24: begin
				q			<=			16'h1793;
		end
		32'h0000AE26: begin
				q			<=			16'h0103;
		end
		32'h0000AE28: begin
				q			<=			16'hD793;
		end
		32'h0000AE2A: begin
				q			<=			16'h0107;
		end
		32'h0000AE2C: begin
				q			<=			16'hE7B3;
		end
		32'h0000AE2E: begin
				q			<=			16'h00F8;
		end
		32'h0000AE30: begin
				q			<=			16'h0713;
		end
		32'h0000AE32: begin
				q			<=			16'h0008;
		end
		32'h0000AE34: begin
				q			<=			16'hFE63;
		end
		32'h0000AE36: begin
				q			<=			16'h01D7;
		end
		32'h0000AE38: begin
				q			<=			16'h87B3;
		end
		32'h0000AE3A: begin
				q			<=			16'h00D7;
		end
		32'h0000AE3C: begin
				q			<=			16'h0713;
		end
		32'h0000AE3E: begin
				q			<=			16'hFFF8;
		end
		32'h0000AE40: begin
				q			<=			16'hE863;
		end
		32'h0000AE42: begin
				q			<=			16'h00D7;
		end
		32'h0000AE44: begin
				q			<=			16'hF663;
		end
		32'h0000AE46: begin
				q			<=			16'h01D7;
		end
		32'h0000AE48: begin
				q			<=			16'h0713;
		end
		32'h0000AE4A: begin
				q			<=			16'hFFE8;
		end
		32'h0000AE4C: begin
				q			<=			16'h87B3;
		end
		32'h0000AE4E: begin
				q			<=			16'h00D7;
		end
		32'h0000AE50: begin
				q			<=			16'h1E13;
		end
		32'h0000AE52: begin
				q			<=			16'h010E;
		end
		32'h0000AE54: begin
				q			<=			16'h87B3;
		end
		32'h0000AE56: begin
				q			<=			16'h41D7;
		end
		32'h0000AE58: begin
				q			<=			16'h0EB7;
		end
		32'h0000AE5A: begin
				q			<=			16'h0001;
		end
		32'h0000AE5C: begin
				q			<=			16'h6733;
		end
		32'h0000AE5E: begin
				q			<=			16'h00EE;
		end
		32'h0000AE60: begin
				q			<=			16'h8813;
		end
		32'h0000AE62: begin
				q			<=			16'hFFFE;
		end
		32'h0000AE64: begin
				q			<=			16'h7333;
		end
		32'h0000AE66: begin
				q			<=			16'h0107;
		end
		32'h0000AE68: begin
				q			<=			16'h5893;
		end
		32'h0000AE6A: begin
				q			<=			16'h0107;
		end
		32'h0000AE6C: begin
				q			<=			16'h7833;
		end
		32'h0000AE6E: begin
				q			<=			16'h0106;
		end
		32'h0000AE70: begin
				q			<=			16'h5613;
		end
		32'h0000AE72: begin
				q			<=			16'h0106;
		end
		32'h0000AE74: begin
				q			<=			16'h0E33;
		end
		32'h0000AE76: begin
				q			<=			16'h0303;
		end
		32'h0000AE78: begin
				q			<=			16'h8833;
		end
		32'h0000AE7A: begin
				q			<=			16'h0308;
		end
		32'h0000AE7C: begin
				q			<=			16'h5693;
		end
		32'h0000AE7E: begin
				q			<=			16'h010E;
		end
		32'h0000AE80: begin
				q			<=			16'h0333;
		end
		32'h0000AE82: begin
				q			<=			16'h02C3;
		end
		32'h0000AE84: begin
				q			<=			16'h0333;
		end
		32'h0000AE86: begin
				q			<=			16'h0103;
		end
		32'h0000AE88: begin
				q			<=			16'h86B3;
		end
		32'h0000AE8A: begin
				q			<=			16'h0066;
		end
		32'h0000AE8C: begin
				q			<=			16'h88B3;
		end
		32'h0000AE8E: begin
				q			<=			16'h02C8;
		end
		32'h0000AE90: begin
				q			<=			16'hF463;
		end
		32'h0000AE92: begin
				q			<=			16'h0106;
		end
		32'h0000AE94: begin
				q			<=			16'h88B3;
		end
		32'h0000AE96: begin
				q			<=			16'h01D8;
		end
		32'h0000AE98: begin
				q			<=			16'hD613;
		end
		32'h0000AE9A: begin
				q			<=			16'h0106;
		end
		32'h0000AE9C: begin
				q			<=			16'h08B3;
		end
		32'h0000AE9E: begin
				q			<=			16'h0116;
		end
		32'h0000AEA0: begin
				q			<=			16'hE663;
		end
		32'h0000AEA2: begin
				q			<=			16'h0317;
		end
		32'h0000AEA4: begin
				q			<=			16'h9AE3;
		end
		32'h0000AEA6: begin
				q			<=			16'hCF17;
		end
		32'h0000AEA8: begin
				q			<=			16'h07B7;
		end
		32'h0000AEAA: begin
				q			<=			16'h0001;
		end
		32'h0000AEAC: begin
				q			<=			16'h8793;
		end
		32'h0000AEAE: begin
				q			<=			16'hFFF7;
		end
		32'h0000AEB0: begin
				q			<=			16'hF6B3;
		end
		32'h0000AEB2: begin
				q			<=			16'h00F6;
		end
		32'h0000AEB4: begin
				q			<=			16'h9693;
		end
		32'h0000AEB6: begin
				q			<=			16'h0106;
		end
		32'h0000AEB8: begin
				q			<=			16'h7E33;
		end
		32'h0000AEBA: begin
				q			<=			16'h00FE;
		end
		32'h0000AEBC: begin
				q			<=			16'h1533;
		end
		32'h0000AEBE: begin
				q			<=			16'h00B5;
		end
		32'h0000AEC0: begin
				q			<=			16'h86B3;
		end
		32'h0000AEC2: begin
				q			<=			16'h01C6;
		end
		32'h0000AEC4: begin
				q			<=			16'h0593;
		end
		32'h0000AEC6: begin
				q			<=			16'h0000;
		end
		32'h0000AEC8: begin
				q			<=			16'h7CE3;
		end
		32'h0000AECA: begin
				q			<=			16'hDAD5;
		end
		32'h0000AECC: begin
				q			<=			16'h0713;
		end
		32'h0000AECE: begin
				q			<=			16'hFFF7;
		end
		32'h0000AED0: begin
				q			<=			16'hF06F;
		end
		32'h0000AED2: begin
				q			<=			16'hCC9F;
		end
		32'h0000AED4: begin
				q			<=			16'h0593;
		end
		32'h0000AED6: begin
				q			<=			16'h0000;
		end
		32'h0000AED8: begin
				q			<=			16'h0713;
		end
		32'h0000AEDA: begin
				q			<=			16'h0000;
		end
		32'h0000AEDC: begin
				q			<=			16'hF06F;
		end
		32'h0000AEDE: begin
				q			<=			16'hDA5F;
		end
		32'h0000AEE0: begin
				q			<=			16'h0000;
		end
		32'h0000AEE2: begin
				q			<=			16'h0000;
		end
		32'h0000AEE4: begin
				q			<=			16'h0893;
		end
		32'h0000AEE6: begin
				q			<=			16'h0006;
		end
		32'h0000AEE8: begin
				q			<=			16'h8713;
		end
		32'h0000AEEA: begin
				q			<=			16'h0006;
		end
		32'h0000AEEC: begin
				q			<=			16'h0793;
		end
		32'h0000AEEE: begin
				q			<=			16'h0005;
		end
		32'h0000AEF0: begin
				q			<=			16'h8813;
		end
		32'h0000AEF2: begin
				q			<=			16'h0005;
		end
		32'h0000AEF4: begin
				q			<=			16'h9C63;
		end
		32'h0000AEF6: begin
				q			<=			16'h2206;
		end
		32'h0000AEF8: begin
				q			<=			16'h5697;
		end
		32'h0000AEFA: begin
				q			<=			16'h0000;
		end
		32'h0000AEFC: begin
				q			<=			16'h8693;
		end
		32'h0000AEFE: begin
				q			<=			16'hA746;
		end
		32'h0000AF00: begin
				q			<=			16'hFC63;
		end
		32'h0000AF02: begin
				q			<=			16'h0CC5;
		end
		32'h0000AF04: begin
				q			<=			16'h0337;
		end
		32'h0000AF06: begin
				q			<=			16'h0001;
		end
		32'h0000AF08: begin
				q			<=			16'h7E63;
		end
		32'h0000AF0A: begin
				q			<=			16'h0A66;
		end
		32'h0000AF0C: begin
				q			<=			16'h0313;
		end
		32'h0000AF0E: begin
				q			<=			16'h0FF0;
		end
		32'h0000AF10: begin
				q			<=			16'h7463;
		end
		32'h0000AF12: begin
				q			<=			16'h00C3;
		end
		32'h0000AF14: begin
				q			<=			16'h0713;
		end
		32'h0000AF16: begin
				q			<=			16'h0080;
		end
		32'h0000AF18: begin
				q			<=			16'h5333;
		end
		32'h0000AF1A: begin
				q			<=			16'h00E6;
		end
		32'h0000AF1C: begin
				q			<=			16'h86B3;
		end
		32'h0000AF1E: begin
				q			<=			16'h0066;
		end
		32'h0000AF20: begin
				q			<=			16'hCE03;
		end
		32'h0000AF22: begin
				q			<=			16'h0006;
		end
		32'h0000AF24: begin
				q			<=			16'h0313;
		end
		32'h0000AF26: begin
				q			<=			16'h0200;
		end
		32'h0000AF28: begin
				q			<=			16'h0E33;
		end
		32'h0000AF2A: begin
				q			<=			16'h00EE;
		end
		32'h0000AF2C: begin
				q			<=			16'h0333;
		end
		32'h0000AF2E: begin
				q			<=			16'h41C3;
		end
		32'h0000AF30: begin
				q			<=			16'h0C63;
		end
		32'h0000AF32: begin
				q			<=			16'h0003;
		end
		32'h0000AF34: begin
				q			<=			16'h95B3;
		end
		32'h0000AF36: begin
				q			<=			16'h0065;
		end
		32'h0000AF38: begin
				q			<=			16'h5E33;
		end
		32'h0000AF3A: begin
				q			<=			16'h01C5;
		end
		32'h0000AF3C: begin
				q			<=			16'h18B3;
		end
		32'h0000AF3E: begin
				q			<=			16'h0066;
		end
		32'h0000AF40: begin
				q			<=			16'h6833;
		end
		32'h0000AF42: begin
				q			<=			16'h00BE;
		end
		32'h0000AF44: begin
				q			<=			16'h17B3;
		end
		32'h0000AF46: begin
				q			<=			16'h0065;
		end
		32'h0000AF48: begin
				q			<=			16'hD613;
		end
		32'h0000AF4A: begin
				q			<=			16'h0108;
		end
		32'h0000AF4C: begin
				q			<=			16'h7733;
		end
		32'h0000AF4E: begin
				q			<=			16'h02C8;
		end
		32'h0000AF50: begin
				q			<=			16'h9513;
		end
		32'h0000AF52: begin
				q			<=			16'h0108;
		end
		32'h0000AF54: begin
				q			<=			16'h5513;
		end
		32'h0000AF56: begin
				q			<=			16'h0105;
		end
		32'h0000AF58: begin
				q			<=			16'hD693;
		end
		32'h0000AF5A: begin
				q			<=			16'h0107;
		end
		32'h0000AF5C: begin
				q			<=			16'h5833;
		end
		32'h0000AF5E: begin
				q			<=			16'h02C8;
		end
		32'h0000AF60: begin
				q			<=			16'h1713;
		end
		32'h0000AF62: begin
				q			<=			16'h0107;
		end
		32'h0000AF64: begin
				q			<=			16'h66B3;
		end
		32'h0000AF66: begin
				q			<=			16'h00D7;
		end
		32'h0000AF68: begin
				q			<=			16'h0833;
		end
		32'h0000AF6A: begin
				q			<=			16'h0305;
		end
		32'h0000AF6C: begin
				q			<=			16'hFA63;
		end
		32'h0000AF6E: begin
				q			<=			16'h0106;
		end
		32'h0000AF70: begin
				q			<=			16'h86B3;
		end
		32'h0000AF72: begin
				q			<=			16'h0116;
		end
		32'h0000AF74: begin
				q			<=			16'hE663;
		end
		32'h0000AF76: begin
				q			<=			16'h0116;
		end
		32'h0000AF78: begin
				q			<=			16'hF463;
		end
		32'h0000AF7A: begin
				q			<=			16'h0106;
		end
		32'h0000AF7C: begin
				q			<=			16'h86B3;
		end
		32'h0000AF7E: begin
				q			<=			16'h0116;
		end
		32'h0000AF80: begin
				q			<=			16'h86B3;
		end
		32'h0000AF82: begin
				q			<=			16'h4106;
		end
		32'h0000AF84: begin
				q			<=			16'hF733;
		end
		32'h0000AF86: begin
				q			<=			16'h02C6;
		end
		32'h0000AF88: begin
				q			<=			16'h9793;
		end
		32'h0000AF8A: begin
				q			<=			16'h0107;
		end
		32'h0000AF8C: begin
				q			<=			16'hD793;
		end
		32'h0000AF8E: begin
				q			<=			16'h0107;
		end
		32'h0000AF90: begin
				q			<=			16'hD6B3;
		end
		32'h0000AF92: begin
				q			<=			16'h02C6;
		end
		32'h0000AF94: begin
				q			<=			16'h06B3;
		end
		32'h0000AF96: begin
				q			<=			16'h02D5;
		end
		32'h0000AF98: begin
				q			<=			16'h1513;
		end
		32'h0000AF9A: begin
				q			<=			16'h0107;
		end
		32'h0000AF9C: begin
				q			<=			16'h67B3;
		end
		32'h0000AF9E: begin
				q			<=			16'h00F5;
		end
		32'h0000AFA0: begin
				q			<=			16'hFA63;
		end
		32'h0000AFA2: begin
				q			<=			16'h00D7;
		end
		32'h0000AFA4: begin
				q			<=			16'h87B3;
		end
		32'h0000AFA6: begin
				q			<=			16'h0117;
		end
		32'h0000AFA8: begin
				q			<=			16'hE663;
		end
		32'h0000AFAA: begin
				q			<=			16'h0117;
		end
		32'h0000AFAC: begin
				q			<=			16'hF463;
		end
		32'h0000AFAE: begin
				q			<=			16'h00D7;
		end
		32'h0000AFB0: begin
				q			<=			16'h87B3;
		end
		32'h0000AFB2: begin
				q			<=			16'h0117;
		end
		32'h0000AFB4: begin
				q			<=			16'h87B3;
		end
		32'h0000AFB6: begin
				q			<=			16'h40D7;
		end
		32'h0000AFB8: begin
				q			<=			16'hD533;
		end
		32'h0000AFBA: begin
				q			<=			16'h0067;
		end
		32'h0000AFBC: begin
				q			<=			16'h0593;
		end
		32'h0000AFBE: begin
				q			<=			16'h0000;
		end
		32'h0000AFC0: begin
				q			<=			16'h8067;
		end
		32'h0000AFC2: begin
				q			<=			16'h0000;
		end
		32'h0000AFC4: begin
				q			<=			16'h0337;
		end
		32'h0000AFC6: begin
				q			<=			16'h0100;
		end
		32'h0000AFC8: begin
				q			<=			16'h0713;
		end
		32'h0000AFCA: begin
				q			<=			16'h0100;
		end
		32'h0000AFCC: begin
				q			<=			16'h66E3;
		end
		32'h0000AFCE: begin
				q			<=			16'hF466;
		end
		32'h0000AFD0: begin
				q			<=			16'h0713;
		end
		32'h0000AFD2: begin
				q			<=			16'h0180;
		end
		32'h0000AFD4: begin
				q			<=			16'hF06F;
		end
		32'h0000AFD6: begin
				q			<=			16'hF45F;
		end
		32'h0000AFD8: begin
				q			<=			16'h1663;
		end
		32'h0000AFDA: begin
				q			<=			16'h0006;
		end
		32'h0000AFDC: begin
				q			<=			16'h0613;
		end
		32'h0000AFDE: begin
				q			<=			16'h0010;
		end
		32'h0000AFE0: begin
				q			<=			16'h58B3;
		end
		32'h0000AFE2: begin
				q			<=			16'h0316;
		end
		32'h0000AFE4: begin
				q			<=			16'h0637;
		end
		32'h0000AFE6: begin
				q			<=			16'h0001;
		end
		32'h0000AFE8: begin
				q			<=			16'hF263;
		end
		32'h0000AFEA: begin
				q			<=			16'h0AC8;
		end
		32'h0000AFEC: begin
				q			<=			16'h0613;
		end
		32'h0000AFEE: begin
				q			<=			16'h0FF0;
		end
		32'h0000AFF0: begin
				q			<=			16'h7463;
		end
		32'h0000AFF2: begin
				q			<=			16'h0116;
		end
		32'h0000AFF4: begin
				q			<=			16'h0713;
		end
		32'h0000AFF6: begin
				q			<=			16'h0080;
		end
		32'h0000AFF8: begin
				q			<=			16'hD633;
		end
		32'h0000AFFA: begin
				q			<=			16'h00E8;
		end
		32'h0000AFFC: begin
				q			<=			16'h86B3;
		end
		32'h0000AFFE: begin
				q			<=			16'h00C6;
		end
		32'h0000B000: begin
				q			<=			16'hCE03;
		end
		32'h0000B002: begin
				q			<=			16'h0006;
		end
		32'h0000B004: begin
				q			<=			16'h0313;
		end
		32'h0000B006: begin
				q			<=			16'h0200;
		end
		32'h0000B008: begin
				q			<=			16'h0E33;
		end
		32'h0000B00A: begin
				q			<=			16'h00EE;
		end
		32'h0000B00C: begin
				q			<=			16'h0333;
		end
		32'h0000B00E: begin
				q			<=			16'h41C3;
		end
		32'h0000B010: begin
				q			<=			16'h1863;
		end
		32'h0000B012: begin
				q			<=			16'h0803;
		end
		32'h0000B014: begin
				q			<=			16'h85B3;
		end
		32'h0000B016: begin
				q			<=			16'h4115;
		end
		32'h0000B018: begin
				q			<=			16'hD713;
		end
		32'h0000B01A: begin
				q			<=			16'h0108;
		end
		32'h0000B01C: begin
				q			<=			16'h9513;
		end
		32'h0000B01E: begin
				q			<=			16'h0108;
		end
		32'h0000B020: begin
				q			<=			16'h5513;
		end
		32'h0000B022: begin
				q			<=			16'h0105;
		end
		32'h0000B024: begin
				q			<=			16'hD613;
		end
		32'h0000B026: begin
				q			<=			16'h0107;
		end
		32'h0000B028: begin
				q			<=			16'hF6B3;
		end
		32'h0000B02A: begin
				q			<=			16'h02E5;
		end
		32'h0000B02C: begin
				q			<=			16'hD5B3;
		end
		32'h0000B02E: begin
				q			<=			16'h02E5;
		end
		32'h0000B030: begin
				q			<=			16'h9693;
		end
		32'h0000B032: begin
				q			<=			16'h0106;
		end
		32'h0000B034: begin
				q			<=			16'hE6B3;
		end
		32'h0000B036: begin
				q			<=			16'h00C6;
		end
		32'h0000B038: begin
				q			<=			16'h05B3;
		end
		32'h0000B03A: begin
				q			<=			16'h02B5;
		end
		32'h0000B03C: begin
				q			<=			16'hFA63;
		end
		32'h0000B03E: begin
				q			<=			16'h00B6;
		end
		32'h0000B040: begin
				q			<=			16'h86B3;
		end
		32'h0000B042: begin
				q			<=			16'h0116;
		end
		32'h0000B044: begin
				q			<=			16'hE663;
		end
		32'h0000B046: begin
				q			<=			16'h0116;
		end
		32'h0000B048: begin
				q			<=			16'hF463;
		end
		32'h0000B04A: begin
				q			<=			16'h00B6;
		end
		32'h0000B04C: begin
				q			<=			16'h86B3;
		end
		32'h0000B04E: begin
				q			<=			16'h0116;
		end
		32'h0000B050: begin
				q			<=			16'h85B3;
		end
		32'h0000B052: begin
				q			<=			16'h40B6;
		end
		32'h0000B054: begin
				q			<=			16'hF6B3;
		end
		32'h0000B056: begin
				q			<=			16'h02E5;
		end
		32'h0000B058: begin
				q			<=			16'h9793;
		end
		32'h0000B05A: begin
				q			<=			16'h0107;
		end
		32'h0000B05C: begin
				q			<=			16'hD793;
		end
		32'h0000B05E: begin
				q			<=			16'h0107;
		end
		32'h0000B060: begin
				q			<=			16'hD5B3;
		end
		32'h0000B062: begin
				q			<=			16'h02E5;
		end
		32'h0000B064: begin
				q			<=			16'h05B3;
		end
		32'h0000B066: begin
				q			<=			16'h02B5;
		end
		32'h0000B068: begin
				q			<=			16'h9513;
		end
		32'h0000B06A: begin
				q			<=			16'h0106;
		end
		32'h0000B06C: begin
				q			<=			16'h67B3;
		end
		32'h0000B06E: begin
				q			<=			16'h00F5;
		end
		32'h0000B070: begin
				q			<=			16'hFA63;
		end
		32'h0000B072: begin
				q			<=			16'h00B7;
		end
		32'h0000B074: begin
				q			<=			16'h87B3;
		end
		32'h0000B076: begin
				q			<=			16'h0117;
		end
		32'h0000B078: begin
				q			<=			16'hE663;
		end
		32'h0000B07A: begin
				q			<=			16'h0117;
		end
		32'h0000B07C: begin
				q			<=			16'hF463;
		end
		32'h0000B07E: begin
				q			<=			16'h00B7;
		end
		32'h0000B080: begin
				q			<=			16'h87B3;
		end
		32'h0000B082: begin
				q			<=			16'h0117;
		end
		32'h0000B084: begin
				q			<=			16'h87B3;
		end
		32'h0000B086: begin
				q			<=			16'h40B7;
		end
		32'h0000B088: begin
				q			<=			16'hF06F;
		end
		32'h0000B08A: begin
				q			<=			16'hF31F;
		end
		32'h0000B08C: begin
				q			<=			16'h0637;
		end
		32'h0000B08E: begin
				q			<=			16'h0100;
		end
		32'h0000B090: begin
				q			<=			16'h0713;
		end
		32'h0000B092: begin
				q			<=			16'h0100;
		end
		32'h0000B094: begin
				q			<=			16'hE2E3;
		end
		32'h0000B096: begin
				q			<=			16'hF6C8;
		end
		32'h0000B098: begin
				q			<=			16'h0713;
		end
		32'h0000B09A: begin
				q			<=			16'h0180;
		end
		32'h0000B09C: begin
				q			<=			16'hF06F;
		end
		32'h0000B09E: begin
				q			<=			16'hF5DF;
		end
		32'h0000B0A0: begin
				q			<=			16'h98B3;
		end
		32'h0000B0A2: begin
				q			<=			16'h0068;
		end
		32'h0000B0A4: begin
				q			<=			16'hD733;
		end
		32'h0000B0A6: begin
				q			<=			16'h01C5;
		end
		32'h0000B0A8: begin
				q			<=			16'h17B3;
		end
		32'h0000B0AA: begin
				q			<=			16'h0065;
		end
		32'h0000B0AC: begin
				q			<=			16'h5E33;
		end
		32'h0000B0AE: begin
				q			<=			16'h01C5;
		end
		32'h0000B0B0: begin
				q			<=			16'hD513;
		end
		32'h0000B0B2: begin
				q			<=			16'h0108;
		end
		32'h0000B0B4: begin
				q			<=			16'h76B3;
		end
		32'h0000B0B6: begin
				q			<=			16'h02A7;
		end
		32'h0000B0B8: begin
				q			<=			16'h95B3;
		end
		32'h0000B0BA: begin
				q			<=			16'h0065;
		end
		32'h0000B0BC: begin
				q			<=			16'h6E33;
		end
		32'h0000B0BE: begin
				q			<=			16'h00BE;
		end
		32'h0000B0C0: begin
				q			<=			16'h9593;
		end
		32'h0000B0C2: begin
				q			<=			16'h0108;
		end
		32'h0000B0C4: begin
				q			<=			16'hD593;
		end
		32'h0000B0C6: begin
				q			<=			16'h0105;
		end
		32'h0000B0C8: begin
				q			<=			16'h5613;
		end
		32'h0000B0CA: begin
				q			<=			16'h010E;
		end
		32'h0000B0CC: begin
				q			<=			16'h5733;
		end
		32'h0000B0CE: begin
				q			<=			16'h02A7;
		end
		32'h0000B0D0: begin
				q			<=			16'h9693;
		end
		32'h0000B0D2: begin
				q			<=			16'h0106;
		end
		32'h0000B0D4: begin
				q			<=			16'hE6B3;
		end
		32'h0000B0D6: begin
				q			<=			16'h00C6;
		end
		32'h0000B0D8: begin
				q			<=			16'h8733;
		end
		32'h0000B0DA: begin
				q			<=			16'h02E5;
		end
		32'h0000B0DC: begin
				q			<=			16'hFA63;
		end
		32'h0000B0DE: begin
				q			<=			16'h00E6;
		end
		32'h0000B0E0: begin
				q			<=			16'h86B3;
		end
		32'h0000B0E2: begin
				q			<=			16'h0116;
		end
		32'h0000B0E4: begin
				q			<=			16'hE663;
		end
		32'h0000B0E6: begin
				q			<=			16'h0116;
		end
		32'h0000B0E8: begin
				q			<=			16'hF463;
		end
		32'h0000B0EA: begin
				q			<=			16'h00E6;
		end
		32'h0000B0EC: begin
				q			<=			16'h86B3;
		end
		32'h0000B0EE: begin
				q			<=			16'h0116;
		end
		32'h0000B0F0: begin
				q			<=			16'h8633;
		end
		32'h0000B0F2: begin
				q			<=			16'h40E6;
		end
		32'h0000B0F4: begin
				q			<=			16'h76B3;
		end
		32'h0000B0F6: begin
				q			<=			16'h02A6;
		end
		32'h0000B0F8: begin
				q			<=			16'h1E13;
		end
		32'h0000B0FA: begin
				q			<=			16'h010E;
		end
		32'h0000B0FC: begin
				q			<=			16'h5E13;
		end
		32'h0000B0FE: begin
				q			<=			16'h010E;
		end
		32'h0000B100: begin
				q			<=			16'h5633;
		end
		32'h0000B102: begin
				q			<=			16'h02A6;
		end
		32'h0000B104: begin
				q			<=			16'h9693;
		end
		32'h0000B106: begin
				q			<=			16'h0106;
		end
		32'h0000B108: begin
				q			<=			16'h8633;
		end
		32'h0000B10A: begin
				q			<=			16'h02C5;
		end
		32'h0000B10C: begin
				q			<=			16'hE5B3;
		end
		32'h0000B10E: begin
				q			<=			16'h01C6;
		end
		32'h0000B110: begin
				q			<=			16'hFA63;
		end
		32'h0000B112: begin
				q			<=			16'h00C5;
		end
		32'h0000B114: begin
				q			<=			16'h85B3;
		end
		32'h0000B116: begin
				q			<=			16'h0115;
		end
		32'h0000B118: begin
				q			<=			16'hE663;
		end
		32'h0000B11A: begin
				q			<=			16'h0115;
		end
		32'h0000B11C: begin
				q			<=			16'hF463;
		end
		32'h0000B11E: begin
				q			<=			16'h00C5;
		end
		32'h0000B120: begin
				q			<=			16'h85B3;
		end
		32'h0000B122: begin
				q			<=			16'h0115;
		end
		32'h0000B124: begin
				q			<=			16'h85B3;
		end
		32'h0000B126: begin
				q			<=			16'h40C5;
		end
		32'h0000B128: begin
				q			<=			16'hF06F;
		end
		32'h0000B12A: begin
				q			<=			16'hEF1F;
		end
		32'h0000B12C: begin
				q			<=			16'hEAE3;
		end
		32'h0000B12E: begin
				q			<=			16'hE8D5;
		end
		32'h0000B130: begin
				q			<=			16'h0737;
		end
		32'h0000B132: begin
				q			<=			16'h0001;
		end
		32'h0000B134: begin
				q			<=			16'hFC63;
		end
		32'h0000B136: begin
				q			<=			16'h04E6;
		end
		32'h0000B138: begin
				q			<=			16'h0E93;
		end
		32'h0000B13A: begin
				q			<=			16'h0FF0;
		end
		32'h0000B13C: begin
				q			<=			16'hB733;
		end
		32'h0000B13E: begin
				q			<=			16'h00DE;
		end
		32'h0000B140: begin
				q			<=			16'h1713;
		end
		32'h0000B142: begin
				q			<=			16'h0037;
		end
		32'h0000B144: begin
				q			<=			16'hD333;
		end
		32'h0000B146: begin
				q			<=			16'h00E6;
		end
		32'h0000B148: begin
				q			<=			16'h5897;
		end
		32'h0000B14A: begin
				q			<=			16'h0000;
		end
		32'h0000B14C: begin
				q			<=			16'h8893;
		end
		32'h0000B14E: begin
				q			<=			16'h8248;
		end
		32'h0000B150: begin
				q			<=			16'h88B3;
		end
		32'h0000B152: begin
				q			<=			16'h0068;
		end
		32'h0000B154: begin
				q			<=			16'hCE83;
		end
		32'h0000B156: begin
				q			<=			16'h0008;
		end
		32'h0000B158: begin
				q			<=			16'h0E13;
		end
		32'h0000B15A: begin
				q			<=			16'h0200;
		end
		32'h0000B15C: begin
				q			<=			16'h8EB3;
		end
		32'h0000B15E: begin
				q			<=			16'h00EE;
		end
		32'h0000B160: begin
				q			<=			16'h0E33;
		end
		32'h0000B162: begin
				q			<=			16'h41DE;
		end
		32'h0000B164: begin
				q			<=			16'h1E63;
		end
		32'h0000B166: begin
				q			<=			16'h020E;
		end
		32'h0000B168: begin
				q			<=			16'hE463;
		end
		32'h0000B16A: begin
				q			<=			16'h00B6;
		end
		32'h0000B16C: begin
				q			<=			16'h6A63;
		end
		32'h0000B16E: begin
				q			<=			16'h00C5;
		end
		32'h0000B170: begin
				q			<=			16'h07B3;
		end
		32'h0000B172: begin
				q			<=			16'h40C5;
		end
		32'h0000B174: begin
				q			<=			16'h85B3;
		end
		32'h0000B176: begin
				q			<=			16'h40D5;
		end
		32'h0000B178: begin
				q			<=			16'h3533;
		end
		32'h0000B17A: begin
				q			<=			16'h00F5;
		end
		32'h0000B17C: begin
				q			<=			16'h8833;
		end
		32'h0000B17E: begin
				q			<=			16'h40A5;
		end
		32'h0000B180: begin
				q			<=			16'h8513;
		end
		32'h0000B182: begin
				q			<=			16'h0007;
		end
		32'h0000B184: begin
				q			<=			16'h0593;
		end
		32'h0000B186: begin
				q			<=			16'h0008;
		end
		32'h0000B188: begin
				q			<=			16'hF06F;
		end
		32'h0000B18A: begin
				q			<=			16'hE39F;
		end
		32'h0000B18C: begin
				q			<=			16'h08B7;
		end
		32'h0000B18E: begin
				q			<=			16'h0100;
		end
		32'h0000B190: begin
				q			<=			16'h0713;
		end
		32'h0000B192: begin
				q			<=			16'h0100;
		end
		32'h0000B194: begin
				q			<=			16'hE8E3;
		end
		32'h0000B196: begin
				q			<=			16'hFB16;
		end
		32'h0000B198: begin
				q			<=			16'h0713;
		end
		32'h0000B19A: begin
				q			<=			16'h0180;
		end
		32'h0000B19C: begin
				q			<=			16'hF06F;
		end
		32'h0000B19E: begin
				q			<=			16'hFA9F;
		end
		32'h0000B1A0: begin
				q			<=			16'h5733;
		end
		32'h0000B1A2: begin
				q			<=			16'h01D6;
		end
		32'h0000B1A4: begin
				q			<=			16'h96B3;
		end
		32'h0000B1A6: begin
				q			<=			16'h01C6;
		end
		32'h0000B1A8: begin
				q			<=			16'h66B3;
		end
		32'h0000B1AA: begin
				q			<=			16'h00D7;
		end
		32'h0000B1AC: begin
				q			<=			16'h57B3;
		end
		32'h0000B1AE: begin
				q			<=			16'h01D5;
		end
		32'h0000B1B0: begin
				q			<=			16'hD733;
		end
		32'h0000B1B2: begin
				q			<=			16'h01D5;
		end
		32'h0000B1B4: begin
				q			<=			16'h95B3;
		end
		32'h0000B1B6: begin
				q			<=			16'h01C5;
		end
		32'h0000B1B8: begin
				q			<=			16'hE7B3;
		end
		32'h0000B1BA: begin
				q			<=			16'h00B7;
		end
		32'h0000B1BC: begin
				q			<=			16'hD593;
		end
		32'h0000B1BE: begin
				q			<=			16'h0106;
		end
		32'h0000B1C0: begin
				q			<=			16'h7333;
		end
		32'h0000B1C2: begin
				q			<=			16'h02B7;
		end
		32'h0000B1C4: begin
				q			<=			16'h9F13;
		end
		32'h0000B1C6: begin
				q			<=			16'h0106;
		end
		32'h0000B1C8: begin
				q			<=			16'h5F13;
		end
		32'h0000B1CA: begin
				q			<=			16'h010F;
		end
		32'h0000B1CC: begin
				q			<=			16'hD893;
		end
		32'h0000B1CE: begin
				q			<=			16'h0107;
		end
		32'h0000B1D0: begin
				q			<=			16'h1633;
		end
		32'h0000B1D2: begin
				q			<=			16'h01C6;
		end
		32'h0000B1D4: begin
				q			<=			16'h1533;
		end
		32'h0000B1D6: begin
				q			<=			16'h01C5;
		end
		32'h0000B1D8: begin
				q			<=			16'h5733;
		end
		32'h0000B1DA: begin
				q			<=			16'h02B7;
		end
		32'h0000B1DC: begin
				q			<=			16'h1313;
		end
		32'h0000B1DE: begin
				q			<=			16'h0103;
		end
		32'h0000B1E0: begin
				q			<=			16'h68B3;
		end
		32'h0000B1E2: begin
				q			<=			16'h0113;
		end
		32'h0000B1E4: begin
				q			<=			16'h0833;
		end
		32'h0000B1E6: begin
				q			<=			16'h02EF;
		end
		32'h0000B1E8: begin
				q			<=			16'h0313;
		end
		32'h0000B1EA: begin
				q			<=			16'h0007;
		end
		32'h0000B1EC: begin
				q			<=			16'hFE63;
		end
		32'h0000B1EE: begin
				q			<=			16'h0108;
		end
		32'h0000B1F0: begin
				q			<=			16'h88B3;
		end
		32'h0000B1F2: begin
				q			<=			16'h00D8;
		end
		32'h0000B1F4: begin
				q			<=			16'h0313;
		end
		32'h0000B1F6: begin
				q			<=			16'hFFF7;
		end
		32'h0000B1F8: begin
				q			<=			16'hE863;
		end
		32'h0000B1FA: begin
				q			<=			16'h00D8;
		end
		32'h0000B1FC: begin
				q			<=			16'hF663;
		end
		32'h0000B1FE: begin
				q			<=			16'h0108;
		end
		32'h0000B200: begin
				q			<=			16'h0313;
		end
		32'h0000B202: begin
				q			<=			16'hFFE7;
		end
		32'h0000B204: begin
				q			<=			16'h88B3;
		end
		32'h0000B206: begin
				q			<=			16'h00D8;
		end
		32'h0000B208: begin
				q			<=			16'h88B3;
		end
		32'h0000B20A: begin
				q			<=			16'h4108;
		end
		32'h0000B20C: begin
				q			<=			16'hFFB3;
		end
		32'h0000B20E: begin
				q			<=			16'h02B8;
		end
		32'h0000B210: begin
				q			<=			16'hD8B3;
		end
		32'h0000B212: begin
				q			<=			16'h02B8;
		end
		32'h0000B214: begin
				q			<=			16'h9F93;
		end
		32'h0000B216: begin
				q			<=			16'h010F;
		end
		32'h0000B218: begin
				q			<=			16'h05B3;
		end
		32'h0000B21A: begin
				q			<=			16'h031F;
		end
		32'h0000B21C: begin
				q			<=			16'h9F13;
		end
		32'h0000B21E: begin
				q			<=			16'h0107;
		end
		32'h0000B220: begin
				q			<=			16'h5F13;
		end
		32'h0000B222: begin
				q			<=			16'h010F;
		end
		32'h0000B224: begin
				q			<=			16'hEF33;
		end
		32'h0000B226: begin
				q			<=			16'h01EF;
		end
		32'h0000B228: begin
				q			<=			16'h8713;
		end
		32'h0000B22A: begin
				q			<=			16'h0008;
		end
		32'h0000B22C: begin
				q			<=			16'h7E63;
		end
		32'h0000B22E: begin
				q			<=			16'h00BF;
		end
		32'h0000B230: begin
				q			<=			16'h0F33;
		end
		32'h0000B232: begin
				q			<=			16'h00DF;
		end
		32'h0000B234: begin
				q			<=			16'h8713;
		end
		32'h0000B236: begin
				q			<=			16'hFFF8;
		end
		32'h0000B238: begin
				q			<=			16'h6863;
		end
		32'h0000B23A: begin
				q			<=			16'h00DF;
		end
		32'h0000B23C: begin
				q			<=			16'h7663;
		end
		32'h0000B23E: begin
				q			<=			16'h00BF;
		end
		32'h0000B240: begin
				q			<=			16'h8713;
		end
		32'h0000B242: begin
				q			<=			16'hFFE8;
		end
		32'h0000B244: begin
				q			<=			16'h0F33;
		end
		32'h0000B246: begin
				q			<=			16'h00DF;
		end
		32'h0000B248: begin
				q			<=			16'h1313;
		end
		32'h0000B24A: begin
				q			<=			16'h0103;
		end
		32'h0000B24C: begin
				q			<=			16'h08B7;
		end
		32'h0000B24E: begin
				q			<=			16'h0001;
		end
		32'h0000B250: begin
				q			<=			16'h6333;
		end
		32'h0000B252: begin
				q			<=			16'h00E3;
		end
		32'h0000B254: begin
				q			<=			16'h8793;
		end
		32'h0000B256: begin
				q			<=			16'hFFF8;
		end
		32'h0000B258: begin
				q			<=			16'h5813;
		end
		32'h0000B25A: begin
				q			<=			16'h0106;
		end
		32'h0000B25C: begin
				q			<=			16'h0F33;
		end
		32'h0000B25E: begin
				q			<=			16'h40BF;
		end
		32'h0000B260: begin
				q			<=			16'h75B3;
		end
		32'h0000B262: begin
				q			<=			16'h00F3;
		end
		32'h0000B264: begin
				q			<=			16'h5313;
		end
		32'h0000B266: begin
				q			<=			16'h0103;
		end
		32'h0000B268: begin
				q			<=			16'h77B3;
		end
		32'h0000B26A: begin
				q			<=			16'h00F6;
		end
		32'h0000B26C: begin
				q			<=			16'h8733;
		end
		32'h0000B26E: begin
				q			<=			16'h02F5;
		end
		32'h0000B270: begin
				q			<=			16'h07B3;
		end
		32'h0000B272: begin
				q			<=			16'h02F3;
		end
		32'h0000B274: begin
				q			<=			16'h85B3;
		end
		32'h0000B276: begin
				q			<=			16'h0305;
		end
		32'h0000B278: begin
				q			<=			16'h0333;
		end
		32'h0000B27A: begin
				q			<=			16'h0303;
		end
		32'h0000B27C: begin
				q			<=			16'h85B3;
		end
		32'h0000B27E: begin
				q			<=			16'h00F5;
		end
		32'h0000B280: begin
				q			<=			16'h5813;
		end
		32'h0000B282: begin
				q			<=			16'h0107;
		end
		32'h0000B284: begin
				q			<=			16'h0833;
		end
		32'h0000B286: begin
				q			<=			16'h00B8;
		end
		32'h0000B288: begin
				q			<=			16'h7463;
		end
		32'h0000B28A: begin
				q			<=			16'h00F8;
		end
		32'h0000B28C: begin
				q			<=			16'h0333;
		end
		32'h0000B28E: begin
				q			<=			16'h0113;
		end
		32'h0000B290: begin
				q			<=			16'h07B7;
		end
		32'h0000B292: begin
				q			<=			16'h0001;
		end
		32'h0000B294: begin
				q			<=			16'h8793;
		end
		32'h0000B296: begin
				q			<=			16'hFFF7;
		end
		32'h0000B298: begin
				q			<=			16'h5593;
		end
		32'h0000B29A: begin
				q			<=			16'h0108;
		end
		32'h0000B29C: begin
				q			<=			16'h7833;
		end
		32'h0000B29E: begin
				q			<=			16'h00F8;
		end
		32'h0000B2A0: begin
				q			<=			16'h1813;
		end
		32'h0000B2A2: begin
				q			<=			16'h0108;
		end
		32'h0000B2A4: begin
				q			<=			16'h7733;
		end
		32'h0000B2A6: begin
				q			<=			16'h00F7;
		end
		32'h0000B2A8: begin
				q			<=			16'h85B3;
		end
		32'h0000B2AA: begin
				q			<=			16'h0065;
		end
		32'h0000B2AC: begin
				q			<=			16'h0733;
		end
		32'h0000B2AE: begin
				q			<=			16'h00E8;
		end
		32'h0000B2B0: begin
				q			<=			16'h6663;
		end
		32'h0000B2B2: begin
				q			<=			16'h00BF;
		end
		32'h0000B2B4: begin
				q			<=			16'h1E63;
		end
		32'h0000B2B6: begin
				q			<=			16'h00BF;
		end
		32'h0000B2B8: begin
				q			<=			16'h7C63;
		end
		32'h0000B2BA: begin
				q			<=			16'h00E5;
		end
		32'h0000B2BC: begin
				q			<=			16'h0633;
		end
		32'h0000B2BE: begin
				q			<=			16'h40C7;
		end
		32'h0000B2C0: begin
				q			<=			16'h3733;
		end
		32'h0000B2C2: begin
				q			<=			16'h00C7;
		end
		32'h0000B2C4: begin
				q			<=			16'h85B3;
		end
		32'h0000B2C6: begin
				q			<=			16'h40D5;
		end
		32'h0000B2C8: begin
				q			<=			16'h85B3;
		end
		32'h0000B2CA: begin
				q			<=			16'h40E5;
		end
		32'h0000B2CC: begin
				q			<=			16'h0713;
		end
		32'h0000B2CE: begin
				q			<=			16'h0006;
		end
		32'h0000B2D0: begin
				q			<=			16'h0733;
		end
		32'h0000B2D2: begin
				q			<=			16'h40E5;
		end
		32'h0000B2D4: begin
				q			<=			16'h3533;
		end
		32'h0000B2D6: begin
				q			<=			16'h00E5;
		end
		32'h0000B2D8: begin
				q			<=			16'h05B3;
		end
		32'h0000B2DA: begin
				q			<=			16'h40BF;
		end
		32'h0000B2DC: begin
				q			<=			16'h85B3;
		end
		32'h0000B2DE: begin
				q			<=			16'h40A5;
		end
		32'h0000B2E0: begin
				q			<=			16'h97B3;
		end
		32'h0000B2E2: begin
				q			<=			16'h01D5;
		end
		32'h0000B2E4: begin
				q			<=			16'h5733;
		end
		32'h0000B2E6: begin
				q			<=			16'h01C7;
		end
		32'h0000B2E8: begin
				q			<=			16'hE533;
		end
		32'h0000B2EA: begin
				q			<=			16'h00E7;
		end
		32'h0000B2EC: begin
				q			<=			16'hD5B3;
		end
		32'h0000B2EE: begin
				q			<=			16'h01C5;
		end
		32'h0000B2F0: begin
				q			<=			16'hF06F;
		end
		32'h0000B2F2: begin
				q			<=			16'hCD1F;
		end
		32'h0000B2F4: begin
				q			<=			16'h0000;
		end
		32'h0000B2F6: begin
				q			<=			16'h0000;
		end
		32'h0000B2F8: begin
				q			<=			16'h0113;
		end
		32'h0000B2FA: begin
				q			<=			16'hFD01;
		end
		32'h0000B2FC: begin
				q			<=			16'h2423;
		end
		32'h0000B2FE: begin
				q			<=			16'h0281;
		end
		32'h0000B300: begin
				q			<=			16'h2223;
		end
		32'h0000B302: begin
				q			<=			16'h0291;
		end
		32'h0000B304: begin
				q			<=			16'h2823;
		end
		32'h0000B306: begin
				q			<=			16'h0161;
		end
		32'h0000B308: begin
				q			<=			16'h0413;
		end
		32'h0000B30A: begin
				q			<=			16'h0005;
		end
		32'h0000B30C: begin
				q			<=			16'h0B13;
		end
		32'h0000B30E: begin
				q			<=			16'h0005;
		end
		32'h0000B310: begin
				q			<=			16'h04B7;
		end
		32'h0000B312: begin
				q			<=			16'h0010;
		end
		32'h0000B314: begin
				q			<=			16'hD513;
		end
		32'h0000B316: begin
				q			<=			16'h0145;
		end
		32'h0000B318: begin
				q			<=			16'h2023;
		end
		32'h0000B31A: begin
				q			<=			16'h0321;
		end
		32'h0000B31C: begin
				q			<=			16'h2E23;
		end
		32'h0000B31E: begin
				q			<=			16'h0131;
		end
		32'h0000B320: begin
				q			<=			16'h2623;
		end
		32'h0000B322: begin
				q			<=			16'h0171;
		end
		32'h0000B324: begin
				q			<=			16'h8493;
		end
		32'h0000B326: begin
				q			<=			16'hFFF4;
		end
		32'h0000B328: begin
				q			<=			16'h2623;
		end
		32'h0000B32A: begin
				q			<=			16'h0211;
		end
		32'h0000B32C: begin
				q			<=			16'h2C23;
		end
		32'h0000B32E: begin
				q			<=			16'h0141;
		end
		32'h0000B330: begin
				q			<=			16'h2A23;
		end
		32'h0000B332: begin
				q			<=			16'h0151;
		end
		32'h0000B334: begin
				q			<=			16'h7513;
		end
		32'h0000B336: begin
				q			<=			16'h7FF5;
		end
		32'h0000B338: begin
				q			<=			16'h0B93;
		end
		32'h0000B33A: begin
				q			<=			16'h0006;
		end
		32'h0000B33C: begin
				q			<=			16'h8993;
		end
		32'h0000B33E: begin
				q			<=			16'h0006;
		end
		32'h0000B340: begin
				q			<=			16'hF4B3;
		end
		32'h0000B342: begin
				q			<=			16'h00B4;
		end
		32'h0000B344: begin
				q			<=			16'hD913;
		end
		32'h0000B346: begin
				q			<=			16'h01F5;
		end
		32'h0000B348: begin
				q			<=			16'h0663;
		end
		32'h0000B34A: begin
				q			<=			16'h0A05;
		end
		32'h0000B34C: begin
				q			<=			16'h0793;
		end
		32'h0000B34E: begin
				q			<=			16'h7FF0;
		end
		32'h0000B350: begin
				q			<=			16'h0663;
		end
		32'h0000B352: begin
				q			<=			16'h10F5;
		end
		32'h0000B354: begin
				q			<=			16'h9493;
		end
		32'h0000B356: begin
				q			<=			16'h0034;
		end
		32'h0000B358: begin
				q			<=			16'h06B7;
		end
		32'h0000B35A: begin
				q			<=			16'h0080;
		end
		32'h0000B35C: begin
				q			<=			16'hE4B3;
		end
		32'h0000B35E: begin
				q			<=			16'h00D4;
		end
		32'h0000B360: begin
				q			<=			16'h5A93;
		end
		32'h0000B362: begin
				q			<=			16'h01DB;
		end
		32'h0000B364: begin
				q			<=			16'hEAB3;
		end
		32'h0000B366: begin
				q			<=			16'h009A;
		end
		32'h0000B368: begin
				q			<=			16'h1413;
		end
		32'h0000B36A: begin
				q			<=			16'h003B;
		end
		32'h0000B36C: begin
				q			<=			16'h0A13;
		end
		32'h0000B36E: begin
				q			<=			16'hC015;
		end
		32'h0000B370: begin
				q			<=			16'h0B13;
		end
		32'h0000B372: begin
				q			<=			16'h0000;
		end
		32'h0000B374: begin
				q			<=			16'hD513;
		end
		32'h0000B376: begin
				q			<=			16'h0149;
		end
		32'h0000B378: begin
				q			<=			16'h04B7;
		end
		32'h0000B37A: begin
				q			<=			16'h0010;
		end
		32'h0000B37C: begin
				q			<=			16'h8493;
		end
		32'h0000B37E: begin
				q			<=			16'hFFF4;
		end
		32'h0000B380: begin
				q			<=			16'h7513;
		end
		32'h0000B382: begin
				q			<=			16'h7FF5;
		end
		32'h0000B384: begin
				q			<=			16'hF4B3;
		end
		32'h0000B386: begin
				q			<=			16'h0134;
		end
		32'h0000B388: begin
				q			<=			16'h8F93;
		end
		32'h0000B38A: begin
				q			<=			16'h000B;
		end
		32'h0000B38C: begin
				q			<=			16'hD993;
		end
		32'h0000B38E: begin
				q			<=			16'h01F9;
		end
		32'h0000B390: begin
				q			<=			16'h0263;
		end
		32'h0000B392: begin
				q			<=			16'h1005;
		end
		32'h0000B394: begin
				q			<=			16'h0793;
		end
		32'h0000B396: begin
				q			<=			16'h7FF0;
		end
		32'h0000B398: begin
				q			<=			16'h0263;
		end
		32'h0000B39A: begin
				q			<=			16'h16F5;
		end
		32'h0000B39C: begin
				q			<=			16'h07B7;
		end
		32'h0000B39E: begin
				q			<=			16'h0080;
		end
		32'h0000B3A0: begin
				q			<=			16'h9493;
		end
		32'h0000B3A2: begin
				q			<=			16'h0034;
		end
		32'h0000B3A4: begin
				q			<=			16'hE4B3;
		end
		32'h0000B3A6: begin
				q			<=			16'h00F4;
		end
		32'h0000B3A8: begin
				q			<=			16'hD793;
		end
		32'h0000B3AA: begin
				q			<=			16'h01DB;
		end
		32'h0000B3AC: begin
				q			<=			16'hE7B3;
		end
		32'h0000B3AE: begin
				q			<=			16'h0097;
		end
		32'h0000B3B0: begin
				q			<=			16'h9F93;
		end
		32'h0000B3B2: begin
				q			<=			16'h003B;
		end
		32'h0000B3B4: begin
				q			<=			16'h0513;
		end
		32'h0000B3B6: begin
				q			<=			16'hC015;
		end
		32'h0000B3B8: begin
				q			<=			16'h0713;
		end
		32'h0000B3BA: begin
				q			<=			16'h0000;
		end
		32'h0000B3BC: begin
				q			<=			16'h1693;
		end
		32'h0000B3BE: begin
				q			<=			16'h002B;
		end
		32'h0000B3C0: begin
				q			<=			16'hE6B3;
		end
		32'h0000B3C2: begin
				q			<=			16'h00E6;
		end
		32'h0000B3C4: begin
				q			<=			16'h8693;
		end
		32'h0000B3C6: begin
				q			<=			16'hFFF6;
		end
		32'h0000B3C8: begin
				q			<=			16'h0593;
		end
		32'h0000B3CA: begin
				q			<=			16'h00E0;
		end
		32'h0000B3CC: begin
				q			<=			16'h4633;
		end
		32'h0000B3CE: begin
				q			<=			16'h0139;
		end
		32'h0000B3D0: begin
				q			<=			16'h0533;
		end
		32'h0000B3D2: begin
				q			<=			16'h40AA;
		end
		32'h0000B3D4: begin
				q			<=			16'hE063;
		end
		32'h0000B3D6: begin
				q			<=			16'h16D5;
		end
		32'h0000B3D8: begin
				q			<=			16'h4597;
		end
		32'h0000B3DA: begin
				q			<=			16'h0000;
		end
		32'h0000B3DC: begin
				q			<=			16'h8593;
		end
		32'h0000B3DE: begin
				q			<=			16'h4E05;
		end
		32'h0000B3E0: begin
				q			<=			16'h9693;
		end
		32'h0000B3E2: begin
				q			<=			16'h0026;
		end
		32'h0000B3E4: begin
				q			<=			16'h86B3;
		end
		32'h0000B3E6: begin
				q			<=			16'h00B6;
		end
		32'h0000B3E8: begin
				q			<=			16'hA683;
		end
		32'h0000B3EA: begin
				q			<=			16'h0006;
		end
		32'h0000B3EC: begin
				q			<=			16'h86B3;
		end
		32'h0000B3EE: begin
				q			<=			16'h00B6;
		end
		32'h0000B3F0: begin
				q			<=			16'h8067;
		end
		32'h0000B3F2: begin
				q			<=			16'h0006;
		end
		32'h0000B3F4: begin
				q			<=			16'hEAB3;
		end
		32'h0000B3F6: begin
				q			<=			16'h0164;
		end
		32'h0000B3F8: begin
				q			<=			16'h8E63;
		end
		32'h0000B3FA: begin
				q			<=			16'h060A;
		end
		32'h0000B3FC: begin
				q			<=			16'h8063;
		end
		32'h0000B3FE: begin
				q			<=			16'h0404;
		end
		32'h0000B400: begin
				q			<=			16'h8513;
		end
		32'h0000B402: begin
				q			<=			16'h0004;
		end
		32'h0000B404: begin
				q			<=			16'h30EF;
		end
		32'h0000B406: begin
				q			<=			16'h4C90;
		end
		32'h0000B408: begin
				q			<=			16'h0793;
		end
		32'h0000B40A: begin
				q			<=			16'hFF55;
		end
		32'h0000B40C: begin
				q			<=			16'h0713;
		end
		32'h0000B40E: begin
				q			<=			16'h01C0;
		end
		32'h0000B410: begin
				q			<=			16'h4E63;
		end
		32'h0000B412: begin
				q			<=			16'h02F7;
		end
		32'h0000B414: begin
				q			<=			16'h0A93;
		end
		32'h0000B416: begin
				q			<=			16'h01D0;
		end
		32'h0000B418: begin
				q			<=			16'h0413;
		end
		32'h0000B41A: begin
				q			<=			16'hFF85;
		end
		32'h0000B41C: begin
				q			<=			16'h8AB3;
		end
		32'h0000B41E: begin
				q			<=			16'h40FA;
		end
		32'h0000B420: begin
				q			<=			16'h94B3;
		end
		32'h0000B422: begin
				q			<=			16'h0084;
		end
		32'h0000B424: begin
				q			<=			16'h5AB3;
		end
		32'h0000B426: begin
				q			<=			16'h015B;
		end
		32'h0000B428: begin
				q			<=			16'hEAB3;
		end
		32'h0000B42A: begin
				q			<=			16'h009A;
		end
		32'h0000B42C: begin
				q			<=			16'h1433;
		end
		32'h0000B42E: begin
				q			<=			16'h008B;
		end
		32'h0000B430: begin
				q			<=			16'h0A13;
		end
		32'h0000B432: begin
				q			<=			16'hC0D0;
		end
		32'h0000B434: begin
				q			<=			16'h0A33;
		end
		32'h0000B436: begin
				q			<=			16'h40AA;
		end
		32'h0000B438: begin
				q			<=			16'hF06F;
		end
		32'h0000B43A: begin
				q			<=			16'hF39F;
		end
		32'h0000B43C: begin
				q			<=			16'h0513;
		end
		32'h0000B43E: begin
				q			<=			16'h000B;
		end
		32'h0000B440: begin
				q			<=			16'h30EF;
		end
		32'h0000B442: begin
				q			<=			16'h48D0;
		end
		32'h0000B444: begin
				q			<=			16'h0513;
		end
		32'h0000B446: begin
				q			<=			16'h0205;
		end
		32'h0000B448: begin
				q			<=			16'hF06F;
		end
		32'h0000B44A: begin
				q			<=			16'hFC1F;
		end
		32'h0000B44C: begin
				q			<=			16'h0493;
		end
		32'h0000B44E: begin
				q			<=			16'hFD85;
		end
		32'h0000B450: begin
				q			<=			16'h1AB3;
		end
		32'h0000B452: begin
				q			<=			16'h009B;
		end
		32'h0000B454: begin
				q			<=			16'h0413;
		end
		32'h0000B456: begin
				q			<=			16'h0000;
		end
		32'h0000B458: begin
				q			<=			16'hF06F;
		end
		32'h0000B45A: begin
				q			<=			16'hFD9F;
		end
		32'h0000B45C: begin
				q			<=			16'hEAB3;
		end
		32'h0000B45E: begin
				q			<=			16'h0164;
		end
		32'h0000B460: begin
				q			<=			16'h8263;
		end
		32'h0000B462: begin
				q			<=			16'h020A;
		end
		32'h0000B464: begin
				q			<=			16'h8A93;
		end
		32'h0000B466: begin
				q			<=			16'h0004;
		end
		32'h0000B468: begin
				q			<=			16'h0A13;
		end
		32'h0000B46A: begin
				q			<=			16'h7FF0;
		end
		32'h0000B46C: begin
				q			<=			16'h0B13;
		end
		32'h0000B46E: begin
				q			<=			16'h0030;
		end
		32'h0000B470: begin
				q			<=			16'hF06F;
		end
		32'h0000B472: begin
				q			<=			16'hF05F;
		end
		32'h0000B474: begin
				q			<=			16'h0413;
		end
		32'h0000B476: begin
				q			<=			16'h0000;
		end
		32'h0000B478: begin
				q			<=			16'h0A13;
		end
		32'h0000B47A: begin
				q			<=			16'h0000;
		end
		32'h0000B47C: begin
				q			<=			16'h0B13;
		end
		32'h0000B47E: begin
				q			<=			16'h0010;
		end
		32'h0000B480: begin
				q			<=			16'hF06F;
		end
		32'h0000B482: begin
				q			<=			16'hEF5F;
		end
		32'h0000B484: begin
				q			<=			16'h0413;
		end
		32'h0000B486: begin
				q			<=			16'h0000;
		end
		32'h0000B488: begin
				q			<=			16'h0A13;
		end
		32'h0000B48A: begin
				q			<=			16'h7FF0;
		end
		32'h0000B48C: begin
				q			<=			16'h0B13;
		end
		32'h0000B48E: begin
				q			<=			16'h0020;
		end
		32'h0000B490: begin
				q			<=			16'hF06F;
		end
		32'h0000B492: begin
				q			<=			16'hEE5F;
		end
		32'h0000B494: begin
				q			<=			16'hE7B3;
		end
		32'h0000B496: begin
				q			<=			16'h0174;
		end
		32'h0000B498: begin
				q			<=			16'h8E63;
		end
		32'h0000B49A: begin
				q			<=			16'h0607;
		end
		32'h0000B49C: begin
				q			<=			16'h8063;
		end
		32'h0000B49E: begin
				q			<=			16'h0404;
		end
		32'h0000B4A0: begin
				q			<=			16'h8513;
		end
		32'h0000B4A2: begin
				q			<=			16'h0004;
		end
		32'h0000B4A4: begin
				q			<=			16'h30EF;
		end
		32'h0000B4A6: begin
				q			<=			16'h4290;
		end
		32'h0000B4A8: begin
				q			<=			16'h0713;
		end
		32'h0000B4AA: begin
				q			<=			16'hFF55;
		end
		32'h0000B4AC: begin
				q			<=			16'h0793;
		end
		32'h0000B4AE: begin
				q			<=			16'h01C0;
		end
		32'h0000B4B0: begin
				q			<=			16'hCE63;
		end
		32'h0000B4B2: begin
				q			<=			16'h02E7;
		end
		32'h0000B4B4: begin
				q			<=			16'h0793;
		end
		32'h0000B4B6: begin
				q			<=			16'h01D0;
		end
		32'h0000B4B8: begin
				q			<=			16'h0F93;
		end
		32'h0000B4BA: begin
				q			<=			16'hFF85;
		end
		32'h0000B4BC: begin
				q			<=			16'h87B3;
		end
		32'h0000B4BE: begin
				q			<=			16'h40E7;
		end
		32'h0000B4C0: begin
				q			<=			16'h94B3;
		end
		32'h0000B4C2: begin
				q			<=			16'h01F4;
		end
		32'h0000B4C4: begin
				q			<=			16'hD7B3;
		end
		32'h0000B4C6: begin
				q			<=			16'h00FB;
		end
		32'h0000B4C8: begin
				q			<=			16'hE7B3;
		end
		32'h0000B4CA: begin
				q			<=			16'h0097;
		end
		32'h0000B4CC: begin
				q			<=			16'h9FB3;
		end
		32'h0000B4CE: begin
				q			<=			16'h01FB;
		end
		32'h0000B4D0: begin
				q			<=			16'h0613;
		end
		32'h0000B4D2: begin
				q			<=			16'hC0D0;
		end
		32'h0000B4D4: begin
				q			<=			16'h0533;
		end
		32'h0000B4D6: begin
				q			<=			16'h40A6;
		end
		32'h0000B4D8: begin
				q			<=			16'hF06F;
		end
		32'h0000B4DA: begin
				q			<=			16'hEE1F;
		end
		32'h0000B4DC: begin
				q			<=			16'h8513;
		end
		32'h0000B4DE: begin
				q			<=			16'h000B;
		end
		32'h0000B4E0: begin
				q			<=			16'h30EF;
		end
		32'h0000B4E2: begin
				q			<=			16'h3ED0;
		end
		32'h0000B4E4: begin
				q			<=			16'h0513;
		end
		32'h0000B4E6: begin
				q			<=			16'h0205;
		end
		32'h0000B4E8: begin
				q			<=			16'hF06F;
		end
		32'h0000B4EA: begin
				q			<=			16'hFC1F;
		end
		32'h0000B4EC: begin
				q			<=			16'h0793;
		end
		32'h0000B4EE: begin
				q			<=			16'hFD85;
		end
		32'h0000B4F0: begin
				q			<=			16'h97B3;
		end
		32'h0000B4F2: begin
				q			<=			16'h00FB;
		end
		32'h0000B4F4: begin
				q			<=			16'h0F93;
		end
		32'h0000B4F6: begin
				q			<=			16'h0000;
		end
		32'h0000B4F8: begin
				q			<=			16'hF06F;
		end
		32'h0000B4FA: begin
				q			<=			16'hFD9F;
		end
		32'h0000B4FC: begin
				q			<=			16'hE7B3;
		end
		32'h0000B4FE: begin
				q			<=			16'h0174;
		end
		32'h0000B500: begin
				q			<=			16'h8263;
		end
		32'h0000B502: begin
				q			<=			16'h0207;
		end
		32'h0000B504: begin
				q			<=			16'h8793;
		end
		32'h0000B506: begin
				q			<=			16'h0004;
		end
		32'h0000B508: begin
				q			<=			16'h0513;
		end
		32'h0000B50A: begin
				q			<=			16'h7FF0;
		end
		32'h0000B50C: begin
				q			<=			16'h0713;
		end
		32'h0000B50E: begin
				q			<=			16'h0030;
		end
		32'h0000B510: begin
				q			<=			16'hF06F;
		end
		32'h0000B512: begin
				q			<=			16'hEADF;
		end
		32'h0000B514: begin
				q			<=			16'h0F93;
		end
		32'h0000B516: begin
				q			<=			16'h0000;
		end
		32'h0000B518: begin
				q			<=			16'h0513;
		end
		32'h0000B51A: begin
				q			<=			16'h0000;
		end
		32'h0000B51C: begin
				q			<=			16'h0713;
		end
		32'h0000B51E: begin
				q			<=			16'h0010;
		end
		32'h0000B520: begin
				q			<=			16'hF06F;
		end
		32'h0000B522: begin
				q			<=			16'hE9DF;
		end
		32'h0000B524: begin
				q			<=			16'h0F93;
		end
		32'h0000B526: begin
				q			<=			16'h0000;
		end
		32'h0000B528: begin
				q			<=			16'h0513;
		end
		32'h0000B52A: begin
				q			<=			16'h7FF0;
		end
		32'h0000B52C: begin
				q			<=			16'h0713;
		end
		32'h0000B52E: begin
				q			<=			16'h0020;
		end
		32'h0000B530: begin
				q			<=			16'hF06F;
		end
		32'h0000B532: begin
				q			<=			16'hE8DF;
		end
		32'h0000B534: begin
				q			<=			16'hE663;
		end
		32'h0000B536: begin
				q			<=			16'h0157;
		end
		32'h0000B538: begin
				q			<=			16'h9063;
		end
		32'h0000B53A: begin
				q			<=			16'h36FA;
		end
		32'h0000B53C: begin
				q			<=			16'h6E63;
		end
		32'h0000B53E: begin
				q			<=			16'h35F4;
		end
		32'h0000B540: begin
				q			<=			16'h9593;
		end
		32'h0000B542: begin
				q			<=			16'h01FA;
		end
		32'h0000B544: begin
				q			<=			16'h5693;
		end
		32'h0000B546: begin
				q			<=			16'h0014;
		end
		32'h0000B548: begin
				q			<=			16'h1713;
		end
		32'h0000B54A: begin
				q			<=			16'h01F4;
		end
		32'h0000B54C: begin
				q			<=			16'hDA93;
		end
		32'h0000B54E: begin
				q			<=			16'h001A;
		end
		32'h0000B550: begin
				q			<=			16'hE433;
		end
		32'h0000B552: begin
				q			<=			16'h00D5;
		end
		32'h0000B554: begin
				q			<=			16'h9793;
		end
		32'h0000B556: begin
				q			<=			16'h0087;
		end
		32'h0000B558: begin
				q			<=			16'hD813;
		end
		32'h0000B55A: begin
				q			<=			16'h018F;
		end
		32'h0000B55C: begin
				q			<=			16'h6833;
		end
		32'h0000B55E: begin
				q			<=			16'h00F8;
		end
		32'h0000B560: begin
				q			<=			16'h5E93;
		end
		32'h0000B562: begin
				q			<=			16'h0108;
		end
		32'h0000B564: begin
				q			<=			16'hD5B3;
		end
		32'h0000B566: begin
				q			<=			16'h03DA;
		end
		32'h0000B568: begin
				q			<=			16'h1E13;
		end
		32'h0000B56A: begin
				q			<=			16'h0108;
		end
		32'h0000B56C: begin
				q			<=			16'h5E13;
		end
		32'h0000B56E: begin
				q			<=			16'h010E;
		end
		32'h0000B570: begin
				q			<=			16'h5693;
		end
		32'h0000B572: begin
				q			<=			16'h0104;
		end
		32'h0000B574: begin
				q			<=			16'h9893;
		end
		32'h0000B576: begin
				q			<=			16'h008F;
		end
		32'h0000B578: begin
				q			<=			16'hF4B3;
		end
		32'h0000B57A: begin
				q			<=			16'h03DA;
		end
		32'h0000B57C: begin
				q			<=			16'h8F93;
		end
		32'h0000B57E: begin
				q			<=			16'h0005;
		end
		32'h0000B580: begin
				q			<=			16'h07B3;
		end
		32'h0000B582: begin
				q			<=			16'h02BE;
		end
		32'h0000B584: begin
				q			<=			16'h9493;
		end
		32'h0000B586: begin
				q			<=			16'h0104;
		end
		32'h0000B588: begin
				q			<=			16'hE6B3;
		end
		32'h0000B58A: begin
				q			<=			16'h0096;
		end
		32'h0000B58C: begin
				q			<=			16'hFE63;
		end
		32'h0000B58E: begin
				q			<=			16'h00F6;
		end
		32'h0000B590: begin
				q			<=			16'h86B3;
		end
		32'h0000B592: begin
				q			<=			16'h0106;
		end
		32'h0000B594: begin
				q			<=			16'h8F93;
		end
		32'h0000B596: begin
				q			<=			16'hFFF5;
		end
		32'h0000B598: begin
				q			<=			16'hE863;
		end
		32'h0000B59A: begin
				q			<=			16'h0106;
		end
		32'h0000B59C: begin
				q			<=			16'hF663;
		end
		32'h0000B59E: begin
				q			<=			16'h00F6;
		end
		32'h0000B5A0: begin
				q			<=			16'h8F93;
		end
		32'h0000B5A2: begin
				q			<=			16'hFFE5;
		end
		32'h0000B5A4: begin
				q			<=			16'h86B3;
		end
		32'h0000B5A6: begin
				q			<=			16'h0106;
		end
		32'h0000B5A8: begin
				q			<=			16'h86B3;
		end
		32'h0000B5AA: begin
				q			<=			16'h40F6;
		end
		32'h0000B5AC: begin
				q			<=			16'hD333;
		end
		32'h0000B5AE: begin
				q			<=			16'h03D6;
		end
		32'h0000B5B0: begin
				q			<=			16'h1413;
		end
		32'h0000B5B2: begin
				q			<=			16'h0104;
		end
		32'h0000B5B4: begin
				q			<=			16'h5413;
		end
		32'h0000B5B6: begin
				q			<=			16'h0104;
		end
		32'h0000B5B8: begin
				q			<=			16'hF6B3;
		end
		32'h0000B5BA: begin
				q			<=			16'h03D6;
		end
		32'h0000B5BC: begin
				q			<=			16'h0793;
		end
		32'h0000B5BE: begin
				q			<=			16'h0003;
		end
		32'h0000B5C0: begin
				q			<=			16'h05B3;
		end
		32'h0000B5C2: begin
				q			<=			16'h026E;
		end
		32'h0000B5C4: begin
				q			<=			16'h9693;
		end
		32'h0000B5C6: begin
				q			<=			16'h0106;
		end
		32'h0000B5C8: begin
				q			<=			16'h66B3;
		end
		32'h0000B5CA: begin
				q			<=			16'h00D4;
		end
		32'h0000B5CC: begin
				q			<=			16'hFE63;
		end
		32'h0000B5CE: begin
				q			<=			16'h00B6;
		end
		32'h0000B5D0: begin
				q			<=			16'h86B3;
		end
		32'h0000B5D2: begin
				q			<=			16'h0106;
		end
		32'h0000B5D4: begin
				q			<=			16'h0793;
		end
		32'h0000B5D6: begin
				q			<=			16'hFFF3;
		end
		32'h0000B5D8: begin
				q			<=			16'hE863;
		end
		32'h0000B5DA: begin
				q			<=			16'h0106;
		end
		32'h0000B5DC: begin
				q			<=			16'hF663;
		end
		32'h0000B5DE: begin
				q			<=			16'h00B6;
		end
		32'h0000B5E0: begin
				q			<=			16'h0793;
		end
		32'h0000B5E2: begin
				q			<=			16'hFFE3;
		end
		32'h0000B5E4: begin
				q			<=			16'h86B3;
		end
		32'h0000B5E6: begin
				q			<=			16'h0106;
		end
		32'h0000B5E8: begin
				q			<=			16'h8433;
		end
		32'h0000B5EA: begin
				q			<=			16'h40B6;
		end
		32'h0000B5EC: begin
				q			<=			16'h9F93;
		end
		32'h0000B5EE: begin
				q			<=			16'h010F;
		end
		32'h0000B5F0: begin
				q			<=			16'h05B7;
		end
		32'h0000B5F2: begin
				q			<=			16'h0001;
		end
		32'h0000B5F4: begin
				q			<=			16'hEFB3;
		end
		32'h0000B5F6: begin
				q			<=			16'h00FF;
		end
		32'h0000B5F8: begin
				q			<=			16'h8313;
		end
		32'h0000B5FA: begin
				q			<=			16'hFFF5;
		end
		32'h0000B5FC: begin
				q			<=			16'hD693;
		end
		32'h0000B5FE: begin
				q			<=			16'h010F;
		end
		32'h0000B600: begin
				q			<=			16'hF7B3;
		end
		32'h0000B602: begin
				q			<=			16'h006F;
		end
		32'h0000B604: begin
				q			<=			16'hDF13;
		end
		32'h0000B606: begin
				q			<=			16'h0108;
		end
		32'h0000B608: begin
				q			<=			16'hF333;
		end
		32'h0000B60A: begin
				q			<=			16'h0068;
		end
		32'h0000B60C: begin
				q			<=			16'h83B3;
		end
		32'h0000B60E: begin
				q			<=			16'h0267;
		end
		32'h0000B610: begin
				q			<=			16'h84B3;
		end
		32'h0000B612: begin
				q			<=			16'h0266;
		end
		32'h0000B614: begin
				q			<=			16'h07B3;
		end
		32'h0000B616: begin
				q			<=			16'h02FF;
		end
		32'h0000B618: begin
				q			<=			16'h82B3;
		end
		32'h0000B61A: begin
				q			<=			16'h03E6;
		end
		32'h0000B61C: begin
				q			<=			16'h86B3;
		end
		32'h0000B61E: begin
				q			<=			16'h0097;
		end
		32'h0000B620: begin
				q			<=			16'hD793;
		end
		32'h0000B622: begin
				q			<=			16'h0103;
		end
		32'h0000B624: begin
				q			<=			16'h87B3;
		end
		32'h0000B626: begin
				q			<=			16'h00D7;
		end
		32'h0000B628: begin
				q			<=			16'hF463;
		end
		32'h0000B62A: begin
				q			<=			16'h0097;
		end
		32'h0000B62C: begin
				q			<=			16'h82B3;
		end
		32'h0000B62E: begin
				q			<=			16'h00B2;
		end
		32'h0000B630: begin
				q			<=			16'hD693;
		end
		32'h0000B632: begin
				q			<=			16'h0107;
		end
		32'h0000B634: begin
				q			<=			16'h86B3;
		end
		32'h0000B636: begin
				q			<=			16'h0056;
		end
		32'h0000B638: begin
				q			<=			16'h02B7;
		end
		32'h0000B63A: begin
				q			<=			16'h0001;
		end
		32'h0000B63C: begin
				q			<=			16'h8293;
		end
		32'h0000B63E: begin
				q			<=			16'hFFF2;
		end
		32'h0000B640: begin
				q			<=			16'hF5B3;
		end
		32'h0000B642: begin
				q			<=			16'h0057;
		end
		32'h0000B644: begin
				q			<=			16'h9593;
		end
		32'h0000B646: begin
				q			<=			16'h0105;
		end
		32'h0000B648: begin
				q			<=			16'hF3B3;
		end
		32'h0000B64A: begin
				q			<=			16'h0053;
		end
		32'h0000B64C: begin
				q			<=			16'h85B3;
		end
		32'h0000B64E: begin
				q			<=			16'h0075;
		end
		32'h0000B650: begin
				q			<=			16'h6863;
		end
		32'h0000B652: begin
				q			<=			16'h00D4;
		end
		32'h0000B654: begin
				q			<=			16'h8793;
		end
		32'h0000B656: begin
				q			<=			16'h000F;
		end
		32'h0000B658: begin
				q			<=			16'h1463;
		end
		32'h0000B65A: begin
				q			<=			16'h04D4;
		end
		32'h0000B65C: begin
				q			<=			16'h7263;
		end
		32'h0000B65E: begin
				q			<=			16'h04B7;
		end
		32'h0000B660: begin
				q			<=			16'h0733;
		end
		32'h0000B662: begin
				q			<=			16'h0117;
		end
		32'h0000B664: begin
				q			<=			16'h32B3;
		end
		32'h0000B666: begin
				q			<=			16'h0117;
		end
		32'h0000B668: begin
				q			<=			16'h82B3;
		end
		32'h0000B66A: begin
				q			<=			16'h0102;
		end
		32'h0000B66C: begin
				q			<=			16'h0433;
		end
		32'h0000B66E: begin
				q			<=			16'h0054;
		end
		32'h0000B670: begin
				q			<=			16'h8793;
		end
		32'h0000B672: begin
				q			<=			16'hFFFF;
		end
		32'h0000B674: begin
				q			<=			16'h6663;
		end
		32'h0000B676: begin
				q			<=			16'h0088;
		end
		32'h0000B678: begin
				q			<=			16'h1463;
		end
		32'h0000B67A: begin
				q			<=			16'h0288;
		end
		32'h0000B67C: begin
				q			<=			16'h6263;
		end
		32'h0000B67E: begin
				q			<=			16'h0317;
		end
		32'h0000B680: begin
				q			<=			16'h6663;
		end
		32'h0000B682: begin
				q			<=			16'h00D4;
		end
		32'h0000B684: begin
				q			<=			16'h9E63;
		end
		32'h0000B686: begin
				q			<=			16'h0086;
		end
		32'h0000B688: begin
				q			<=			16'h7C63;
		end
		32'h0000B68A: begin
				q			<=			16'h00B7;
		end
		32'h0000B68C: begin
				q			<=			16'h0733;
		end
		32'h0000B68E: begin
				q			<=			16'h0117;
		end
		32'h0000B690: begin
				q			<=			16'h8793;
		end
		32'h0000B692: begin
				q			<=			16'hFFEF;
		end
		32'h0000B694: begin
				q			<=			16'h3FB3;
		end
		32'h0000B696: begin
				q			<=			16'h0117;
		end
		32'h0000B698: begin
				q			<=			16'h8FB3;
		end
		32'h0000B69A: begin
				q			<=			16'h010F;
		end
		32'h0000B69C: begin
				q			<=			16'h0433;
		end
		32'h0000B69E: begin
				q			<=			16'h01F4;
		end
		32'h0000B6A0: begin
				q			<=			16'h05B3;
		end
		32'h0000B6A2: begin
				q			<=			16'h40B7;
		end
		32'h0000B6A4: begin
				q			<=			16'h0433;
		end
		32'h0000B6A6: begin
				q			<=			16'h40D4;
		end
		32'h0000B6A8: begin
				q			<=			16'h3733;
		end
		32'h0000B6AA: begin
				q			<=			16'h00B7;
		end
		32'h0000B6AC: begin
				q			<=			16'h0433;
		end
		32'h0000B6AE: begin
				q			<=			16'h40E4;
		end
		32'h0000B6B0: begin
				q			<=			16'h0F93;
		end
		32'h0000B6B2: begin
				q			<=			16'hFFF0;
		end
		32'h0000B6B4: begin
				q			<=			16'h0463;
		end
		32'h0000B6B6: begin
				q			<=			16'h1288;
		end
		32'h0000B6B8: begin
				q			<=			16'h52B3;
		end
		32'h0000B6BA: begin
				q			<=			16'h03D4;
		end
		32'h0000B6BC: begin
				q			<=			16'hD693;
		end
		32'h0000B6BE: begin
				q			<=			16'h0105;
		end
		32'h0000B6C0: begin
				q			<=			16'h7433;
		end
		32'h0000B6C2: begin
				q			<=			16'h03D4;
		end
		32'h0000B6C4: begin
				q			<=			16'h8713;
		end
		32'h0000B6C6: begin
				q			<=			16'h0002;
		end
		32'h0000B6C8: begin
				q			<=			16'h0FB3;
		end
		32'h0000B6CA: begin
				q			<=			16'h025E;
		end
		32'h0000B6CC: begin
				q			<=			16'h1413;
		end
		32'h0000B6CE: begin
				q			<=			16'h0104;
		end
		32'h0000B6D0: begin
				q			<=			16'hE433;
		end
		32'h0000B6D2: begin
				q			<=			16'h0086;
		end
		32'h0000B6D4: begin
				q			<=			16'h7E63;
		end
		32'h0000B6D6: begin
				q			<=			16'h01F4;
		end
		32'h0000B6D8: begin
				q			<=			16'h0433;
		end
		32'h0000B6DA: begin
				q			<=			16'h0104;
		end
		32'h0000B6DC: begin
				q			<=			16'h8713;
		end
		32'h0000B6DE: begin
				q			<=			16'hFFF2;
		end
		32'h0000B6E0: begin
				q			<=			16'h6863;
		end
		32'h0000B6E2: begin
				q			<=			16'h0104;
		end
		32'h0000B6E4: begin
				q			<=			16'h7663;
		end
		32'h0000B6E6: begin
				q			<=			16'h01F4;
		end
		32'h0000B6E8: begin
				q			<=			16'h8713;
		end
		32'h0000B6EA: begin
				q			<=			16'hFFE2;
		end
		32'h0000B6EC: begin
				q			<=			16'h0433;
		end
		32'h0000B6EE: begin
				q			<=			16'h0104;
		end
		32'h0000B6F0: begin
				q			<=			16'h0433;
		end
		32'h0000B6F2: begin
				q			<=			16'h41F4;
		end
		32'h0000B6F4: begin
				q			<=			16'h56B3;
		end
		32'h0000B6F6: begin
				q			<=			16'h03D4;
		end
		32'h0000B6F8: begin
				q			<=			16'h9593;
		end
		32'h0000B6FA: begin
				q			<=			16'h0105;
		end
		32'h0000B6FC: begin
				q			<=			16'hD593;
		end
		32'h0000B6FE: begin
				q			<=			16'h0105;
		end
		32'h0000B700: begin
				q			<=			16'h7433;
		end
		32'h0000B702: begin
				q			<=			16'h03D4;
		end
		32'h0000B704: begin
				q			<=			16'h0E33;
		end
		32'h0000B706: begin
				q			<=			16'h02DE;
		end
		32'h0000B708: begin
				q			<=			16'h1413;
		end
		32'h0000B70A: begin
				q			<=			16'h0104;
		end
		32'h0000B70C: begin
				q			<=			16'hE433;
		end
		32'h0000B70E: begin
				q			<=			16'h0085;
		end
		32'h0000B710: begin
				q			<=			16'h8593;
		end
		32'h0000B712: begin
				q			<=			16'h0006;
		end
		32'h0000B714: begin
				q			<=			16'h7E63;
		end
		32'h0000B716: begin
				q			<=			16'h01C4;
		end
		32'h0000B718: begin
				q			<=			16'h0433;
		end
		32'h0000B71A: begin
				q			<=			16'h0104;
		end
		32'h0000B71C: begin
				q			<=			16'h8593;
		end
		32'h0000B71E: begin
				q			<=			16'hFFF6;
		end
		32'h0000B720: begin
				q			<=			16'h6863;
		end
		32'h0000B722: begin
				q			<=			16'h0104;
		end
		32'h0000B724: begin
				q			<=			16'h7663;
		end
		32'h0000B726: begin
				q			<=			16'h01C4;
		end
		32'h0000B728: begin
				q			<=			16'h8593;
		end
		32'h0000B72A: begin
				q			<=			16'hFFE6;
		end
		32'h0000B72C: begin
				q			<=			16'h0433;
		end
		32'h0000B72E: begin
				q			<=			16'h0104;
		end
		32'h0000B730: begin
				q			<=			16'h1713;
		end
		32'h0000B732: begin
				q			<=			16'h0107;
		end
		32'h0000B734: begin
				q			<=			16'h65B3;
		end
		32'h0000B736: begin
				q			<=			16'h00B7;
		end
		32'h0000B738: begin
				q			<=			16'h9713;
		end
		32'h0000B73A: begin
				q			<=			16'h0105;
		end
		32'h0000B73C: begin
				q			<=			16'h5713;
		end
		32'h0000B73E: begin
				q			<=			16'h0107;
		end
		32'h0000B740: begin
				q			<=			16'h0433;
		end
		32'h0000B742: begin
				q			<=			16'h41C4;
		end
		32'h0000B744: begin
				q			<=			16'hDE13;
		end
		32'h0000B746: begin
				q			<=			16'h0105;
		end
		32'h0000B748: begin
				q			<=			16'h0EB3;
		end
		32'h0000B74A: begin
				q			<=			16'h0267;
		end
		32'h0000B74C: begin
				q			<=			16'h0333;
		end
		32'h0000B74E: begin
				q			<=			16'h026E;
		end
		32'h0000B750: begin
				q			<=			16'h0E33;
		end
		32'h0000B752: begin
				q			<=			16'h03CF;
		end
		32'h0000B754: begin
				q			<=			16'h0F33;
		end
		32'h0000B756: begin
				q			<=			16'h02EF;
		end
		32'h0000B758: begin
				q			<=			16'hD713;
		end
		32'h0000B75A: begin
				q			<=			16'h010E;
		end
		32'h0000B75C: begin
				q			<=			16'h0F33;
		end
		32'h0000B75E: begin
				q			<=			16'h006F;
		end
		32'h0000B760: begin
				q			<=			16'h0733;
		end
		32'h0000B762: begin
				q			<=			16'h01E7;
		end
		32'h0000B764: begin
				q			<=			16'h7663;
		end
		32'h0000B766: begin
				q			<=			16'h0067;
		end
		32'h0000B768: begin
				q			<=			16'h06B7;
		end
		32'h0000B76A: begin
				q			<=			16'h0001;
		end
		32'h0000B76C: begin
				q			<=			16'h0E33;
		end
		32'h0000B76E: begin
				q			<=			16'h00DE;
		end
		32'h0000B770: begin
				q			<=			16'h5313;
		end
		32'h0000B772: begin
				q			<=			16'h0107;
		end
		32'h0000B774: begin
				q			<=			16'h0333;
		end
		32'h0000B776: begin
				q			<=			16'h01C3;
		end
		32'h0000B778: begin
				q			<=			16'h0E37;
		end
		32'h0000B77A: begin
				q			<=			16'h0001;
		end
		32'h0000B77C: begin
				q			<=			16'h0E13;
		end
		32'h0000B77E: begin
				q			<=			16'hFFFE;
		end
		32'h0000B780: begin
				q			<=			16'h76B3;
		end
		32'h0000B782: begin
				q			<=			16'h01C7;
		end
		32'h0000B784: begin
				q			<=			16'h9693;
		end
		32'h0000B786: begin
				q			<=			16'h0106;
		end
		32'h0000B788: begin
				q			<=			16'hFEB3;
		end
		32'h0000B78A: begin
				q			<=			16'h01CE;
		end
		32'h0000B78C: begin
				q			<=			16'h86B3;
		end
		32'h0000B78E: begin
				q			<=			16'h01D6;
		end
		32'h0000B790: begin
				q			<=			16'h6863;
		end
		32'h0000B792: begin
				q			<=			16'h0064;
		end
		32'h0000B794: begin
				q			<=			16'h8F93;
		end
		32'h0000B796: begin
				q			<=			16'h0005;
		end
		32'h0000B798: begin
				q			<=			16'h1063;
		end
		32'h0000B79A: begin
				q			<=			16'h0464;
		end
		32'h0000B79C: begin
				q			<=			16'h8063;
		end
		32'h0000B79E: begin
				q			<=			16'h0406;
		end
		32'h0000B7A0: begin
				q			<=			16'h0433;
		end
		32'h0000B7A2: begin
				q			<=			16'h0088;
		end
		32'h0000B7A4: begin
				q			<=			16'h8F93;
		end
		32'h0000B7A6: begin
				q			<=			16'hFFF5;
		end
		32'h0000B7A8: begin
				q			<=			16'h6463;
		end
		32'h0000B7AA: begin
				q			<=			16'h0304;
		end
		32'h0000B7AC: begin
				q			<=			16'h6663;
		end
		32'h0000B7AE: begin
				q			<=			16'h0064;
		end
		32'h0000B7B0: begin
				q			<=			16'h1463;
		end
		32'h0000B7B2: begin
				q			<=			16'h0264;
		end
		32'h0000B7B4: begin
				q			<=			16'hF063;
		end
		32'h0000B7B6: begin
				q			<=			16'h02D8;
		end
		32'h0000B7B8: begin
				q			<=			16'h9713;
		end
		32'h0000B7BA: begin
				q			<=			16'h0018;
		end
		32'h0000B7BC: begin
				q			<=			16'h38B3;
		end
		32'h0000B7BE: begin
				q			<=			16'h0117;
		end
		32'h0000B7C0: begin
				q			<=			16'h8833;
		end
		32'h0000B7C2: begin
				q			<=			16'h0108;
		end
		32'h0000B7C4: begin
				q			<=			16'h8F93;
		end
		32'h0000B7C6: begin
				q			<=			16'hFFE5;
		end
		32'h0000B7C8: begin
				q			<=			16'h0433;
		end
		32'h0000B7CA: begin
				q			<=			16'h0104;
		end
		32'h0000B7CC: begin
				q			<=			16'h0893;
		end
		32'h0000B7CE: begin
				q			<=			16'h0007;
		end
		32'h0000B7D0: begin
				q			<=			16'h1463;
		end
		32'h0000B7D2: begin
				q			<=			16'h0064;
		end
		32'h0000B7D4: begin
				q			<=			16'h8463;
		end
		32'h0000B7D6: begin
				q			<=			16'h0116;
		end
		32'h0000B7D8: begin
				q			<=			16'hEF93;
		end
		32'h0000B7DA: begin
				q			<=			16'h001F;
		end
		32'h0000B7DC: begin
				q			<=			16'h0693;
		end
		32'h0000B7DE: begin
				q			<=			16'h3FF5;
		end
		32'h0000B7E0: begin
				q			<=			16'h5A63;
		end
		32'h0000B7E2: begin
				q			<=			16'h10D0;
		end
		32'h0000B7E4: begin
				q			<=			16'hF713;
		end
		32'h0000B7E6: begin
				q			<=			16'h007F;
		end
		32'h0000B7E8: begin
				q			<=			16'h0063;
		end
		32'h0000B7EA: begin
				q			<=			16'h0207;
		end
		32'h0000B7EC: begin
				q			<=			16'hF713;
		end
		32'h0000B7EE: begin
				q			<=			16'h00FF;
		end
		32'h0000B7F0: begin
				q			<=			16'h0593;
		end
		32'h0000B7F2: begin
				q			<=			16'h0040;
		end
		32'h0000B7F4: begin
				q			<=			16'h0A63;
		end
		32'h0000B7F6: begin
				q			<=			16'h00B7;
		end
		32'h0000B7F8: begin
				q			<=			16'h8593;
		end
		32'h0000B7FA: begin
				q			<=			16'h004F;
		end
		32'h0000B7FC: begin
				q			<=			16'hBFB3;
		end
		32'h0000B7FE: begin
				q			<=			16'h01F5;
		end
		32'h0000B800: begin
				q			<=			16'h87B3;
		end
		32'h0000B802: begin
				q			<=			16'h01F7;
		end
		32'h0000B804: begin
				q			<=			16'h8F93;
		end
		32'h0000B806: begin
				q			<=			16'h0005;
		end
		32'h0000B808: begin
				q			<=			16'h9713;
		end
		32'h0000B80A: begin
				q			<=			16'h0077;
		end
		32'h0000B80C: begin
				q			<=			16'h5A63;
		end
		32'h0000B80E: begin
				q			<=			16'h0007;
		end
		32'h0000B810: begin
				q			<=			16'h0737;
		end
		32'h0000B812: begin
				q			<=			16'hFF00;
		end
		32'h0000B814: begin
				q			<=			16'h0713;
		end
		32'h0000B816: begin
				q			<=			16'hFFF7;
		end
		32'h0000B818: begin
				q			<=			16'hF7B3;
		end
		32'h0000B81A: begin
				q			<=			16'h00E7;
		end
		32'h0000B81C: begin
				q			<=			16'h0693;
		end
		32'h0000B81E: begin
				q			<=			16'h4005;
		end
		32'h0000B820: begin
				q			<=			16'h0713;
		end
		32'h0000B822: begin
				q			<=			16'h7FE0;
		end
		32'h0000B824: begin
				q			<=			16'h4A63;
		end
		32'h0000B826: begin
				q			<=			16'h18D7;
		end
		32'h0000B828: begin
				q			<=			16'h9713;
		end
		32'h0000B82A: begin
				q			<=			16'h01D7;
		end
		32'h0000B82C: begin
				q			<=			16'hDF93;
		end
		32'h0000B82E: begin
				q			<=			16'h003F;
		end
		32'h0000B830: begin
				q			<=			16'h6733;
		end
		32'h0000B832: begin
				q			<=			16'h01F7;
		end
		32'h0000B834: begin
				q			<=			16'hD793;
		end
		32'h0000B836: begin
				q			<=			16'h0037;
		end
		32'h0000B838: begin
				q			<=			16'h05B7;
		end
		32'h0000B83A: begin
				q			<=			16'h0010;
		end
		32'h0000B83C: begin
				q			<=			16'h8593;
		end
		32'h0000B83E: begin
				q			<=			16'hFFF5;
		end
		32'h0000B840: begin
				q			<=			16'hF7B3;
		end
		32'h0000B842: begin
				q			<=			16'h00B7;
		end
		32'h0000B844: begin
				q			<=			16'h05B7;
		end
		32'h0000B846: begin
				q			<=			16'h8010;
		end
		32'h0000B848: begin
				q			<=			16'h8593;
		end
		32'h0000B84A: begin
				q			<=			16'hFFF5;
		end
		32'h0000B84C: begin
				q			<=			16'hF693;
		end
		32'h0000B84E: begin
				q			<=			16'h7FF6;
		end
		32'h0000B850: begin
				q			<=			16'h9693;
		end
		32'h0000B852: begin
				q			<=			16'h0146;
		end
		32'h0000B854: begin
				q			<=			16'hF7B3;
		end
		32'h0000B856: begin
				q			<=			16'h00B7;
		end
		32'h0000B858: begin
				q			<=			16'h2083;
		end
		32'h0000B85A: begin
				q			<=			16'h02C1;
		end
		32'h0000B85C: begin
				q			<=			16'h2403;
		end
		32'h0000B85E: begin
				q			<=			16'h0281;
		end
		32'h0000B860: begin
				q			<=			16'h1613;
		end
		32'h0000B862: begin
				q			<=			16'h01F6;
		end
		32'h0000B864: begin
				q			<=			16'hE7B3;
		end
		32'h0000B866: begin
				q			<=			16'h00D7;
		end
		32'h0000B868: begin
				q			<=			16'hE6B3;
		end
		32'h0000B86A: begin
				q			<=			16'h00C7;
		end
		32'h0000B86C: begin
				q			<=			16'h2483;
		end
		32'h0000B86E: begin
				q			<=			16'h0241;
		end
		32'h0000B870: begin
				q			<=			16'h2903;
		end
		32'h0000B872: begin
				q			<=			16'h0201;
		end
		32'h0000B874: begin
				q			<=			16'h2983;
		end
		32'h0000B876: begin
				q			<=			16'h01C1;
		end
		32'h0000B878: begin
				q			<=			16'h2A03;
		end
		32'h0000B87A: begin
				q			<=			16'h0181;
		end
		32'h0000B87C: begin
				q			<=			16'h2A83;
		end
		32'h0000B87E: begin
				q			<=			16'h0141;
		end
		32'h0000B880: begin
				q			<=			16'h2B03;
		end
		32'h0000B882: begin
				q			<=			16'h0101;
		end
		32'h0000B884: begin
				q			<=			16'h2B83;
		end
		32'h0000B886: begin
				q			<=			16'h00C1;
		end
		32'h0000B888: begin
				q			<=			16'h0513;
		end
		32'h0000B88A: begin
				q			<=			16'h0007;
		end
		32'h0000B88C: begin
				q			<=			16'h8593;
		end
		32'h0000B88E: begin
				q			<=			16'h0006;
		end
		32'h0000B890: begin
				q			<=			16'h0113;
		end
		32'h0000B892: begin
				q			<=			16'h0301;
		end
		32'h0000B894: begin
				q			<=			16'h8067;
		end
		32'h0000B896: begin
				q			<=			16'h0000;
		end
		32'h0000B898: begin
				q			<=			16'h0513;
		end
		32'h0000B89A: begin
				q			<=			16'hFFF5;
		end
		32'h0000B89C: begin
				q			<=			16'h0713;
		end
		32'h0000B89E: begin
				q			<=			16'h0000;
		end
		32'h0000B8A0: begin
				q			<=			16'hF06F;
		end
		32'h0000B8A2: begin
				q			<=			16'hCB5F;
		end
		32'h0000B8A4: begin
				q			<=			16'h0613;
		end
		32'h0000B8A6: begin
				q			<=			16'h0009;
		end
		32'h0000B8A8: begin
				q			<=			16'h8793;
		end
		32'h0000B8AA: begin
				q			<=			16'h000A;
		end
		32'h0000B8AC: begin
				q			<=			16'h0F93;
		end
		32'h0000B8AE: begin
				q			<=			16'h0004;
		end
		32'h0000B8B0: begin
				q			<=			16'h0713;
		end
		32'h0000B8B2: begin
				q			<=			16'h000B;
		end
		32'h0000B8B4: begin
				q			<=			16'h0693;
		end
		32'h0000B8B6: begin
				q			<=			16'h0020;
		end
		32'h0000B8B8: begin
				q			<=			16'h0063;
		end
		32'h0000B8BA: begin
				q			<=			16'h10D7;
		end
		32'h0000B8BC: begin
				q			<=			16'h0693;
		end
		32'h0000B8BE: begin
				q			<=			16'h0030;
		end
		32'h0000B8C0: begin
				q			<=			16'h0263;
		end
		32'h0000B8C2: begin
				q			<=			16'h0ED7;
		end
		32'h0000B8C4: begin
				q			<=			16'h0693;
		end
		32'h0000B8C6: begin
				q			<=			16'h0010;
		end
		32'h0000B8C8: begin
				q			<=			16'h1AE3;
		end
		32'h0000B8CA: begin
				q			<=			16'hF0D7;
		end
		32'h0000B8CC: begin
				q			<=			16'h0793;
		end
		32'h0000B8CE: begin
				q			<=			16'h0000;
		end
		32'h0000B8D0: begin
				q			<=			16'h0713;
		end
		32'h0000B8D2: begin
				q			<=			16'h0000;
		end
		32'h0000B8D4: begin
				q			<=			16'h006F;
		end
		32'h0000B8D6: begin
				q			<=			16'h0940;
		end
		32'h0000B8D8: begin
				q			<=			16'h8613;
		end
		32'h0000B8DA: begin
				q			<=			16'h0009;
		end
		32'h0000B8DC: begin
				q			<=			16'hF06F;
		end
		32'h0000B8DE: begin
				q			<=			16'hFD9F;
		end
		32'h0000B8E0: begin
				q			<=			16'h07B7;
		end
		32'h0000B8E2: begin
				q			<=			16'h0008;
		end
		32'h0000B8E4: begin
				q			<=			16'h0F93;
		end
		32'h0000B8E6: begin
				q			<=			16'h0000;
		end
		32'h0000B8E8: begin
				q			<=			16'h0613;
		end
		32'h0000B8EA: begin
				q			<=			16'h0000;
		end
		32'h0000B8EC: begin
				q			<=			16'h0713;
		end
		32'h0000B8EE: begin
				q			<=			16'h0030;
		end
		32'h0000B8F0: begin
				q			<=			16'hF06F;
		end
		32'h0000B8F2: begin
				q			<=			16'hFC5F;
		end
		32'h0000B8F4: begin
				q			<=			16'h0593;
		end
		32'h0000B8F6: begin
				q			<=			16'h0010;
		end
		32'h0000B8F8: begin
				q			<=			16'h85B3;
		end
		32'h0000B8FA: begin
				q			<=			16'h40D5;
		end
		32'h0000B8FC: begin
				q			<=			16'h0713;
		end
		32'h0000B8FE: begin
				q			<=			16'h0380;
		end
		32'h0000B900: begin
				q			<=			16'h46E3;
		end
		32'h0000B902: begin
				q			<=			16'hFCB7;
		end
		32'h0000B904: begin
				q			<=			16'h0713;
		end
		32'h0000B906: begin
				q			<=			16'h01F0;
		end
		32'h0000B908: begin
				q			<=			16'h4463;
		end
		32'h0000B90A: begin
				q			<=			16'h06B7;
		end
		32'h0000B90C: begin
				q			<=			16'h0513;
		end
		32'h0000B90E: begin
				q			<=			16'h41E5;
		end
		32'h0000B910: begin
				q			<=			16'h9733;
		end
		32'h0000B912: begin
				q			<=			16'h00A7;
		end
		32'h0000B914: begin
				q			<=			16'hD6B3;
		end
		32'h0000B916: begin
				q			<=			16'h00BF;
		end
		32'h0000B918: begin
				q			<=			16'h9533;
		end
		32'h0000B91A: begin
				q			<=			16'h00AF;
		end
		32'h0000B91C: begin
				q			<=			16'h6733;
		end
		32'h0000B91E: begin
				q			<=			16'h00D7;
		end
		32'h0000B920: begin
				q			<=			16'h3533;
		end
		32'h0000B922: begin
				q			<=			16'h00A0;
		end
		32'h0000B924: begin
				q			<=			16'h6733;
		end
		32'h0000B926: begin
				q			<=			16'h00A7;
		end
		32'h0000B928: begin
				q			<=			16'hD7B3;
		end
		32'h0000B92A: begin
				q			<=			16'h00B7;
		end
		32'h0000B92C: begin
				q			<=			16'h7693;
		end
		32'h0000B92E: begin
				q			<=			16'h0077;
		end
		32'h0000B930: begin
				q			<=			16'h8063;
		end
		32'h0000B932: begin
				q			<=			16'h0206;
		end
		32'h0000B934: begin
				q			<=			16'h7693;
		end
		32'h0000B936: begin
				q			<=			16'h00F7;
		end
		32'h0000B938: begin
				q			<=			16'h0593;
		end
		32'h0000B93A: begin
				q			<=			16'h0040;
		end
		32'h0000B93C: begin
				q			<=			16'h8A63;
		end
		32'h0000B93E: begin
				q			<=			16'h00B6;
		end
		32'h0000B940: begin
				q			<=			16'h0693;
		end
		32'h0000B942: begin
				q			<=			16'h0047;
		end
		32'h0000B944: begin
				q			<=			16'hB733;
		end
		32'h0000B946: begin
				q			<=			16'h00E6;
		end
		32'h0000B948: begin
				q			<=			16'h87B3;
		end
		32'h0000B94A: begin
				q			<=			16'h00E7;
		end
		32'h0000B94C: begin
				q			<=			16'h8713;
		end
		32'h0000B94E: begin
				q			<=			16'h0006;
		end
		32'h0000B950: begin
				q			<=			16'h9693;
		end
		32'h0000B952: begin
				q			<=			16'h0087;
		end
		32'h0000B954: begin
				q			<=			16'hCA63;
		end
		32'h0000B956: begin
				q			<=			16'h0606;
		end
		32'h0000B958: begin
				q			<=			16'h9693;
		end
		32'h0000B95A: begin
				q			<=			16'h01D7;
		end
		32'h0000B95C: begin
				q			<=			16'h5713;
		end
		32'h0000B95E: begin
				q			<=			16'h0037;
		end
		32'h0000B960: begin
				q			<=			16'hE733;
		end
		32'h0000B962: begin
				q			<=			16'h00E6;
		end
		32'h0000B964: begin
				q			<=			16'hD793;
		end
		32'h0000B966: begin
				q			<=			16'h0037;
		end
		32'h0000B968: begin
				q			<=			16'h0693;
		end
		32'h0000B96A: begin
				q			<=			16'h0000;
		end
		32'h0000B96C: begin
				q			<=			16'hF06F;
		end
		32'h0000B96E: begin
				q			<=			16'hECDF;
		end
		32'h0000B970: begin
				q			<=			16'h0713;
		end
		32'h0000B972: begin
				q			<=			16'hFE10;
		end
		32'h0000B974: begin
				q			<=			16'h0733;
		end
		32'h0000B976: begin
				q			<=			16'h40D7;
		end
		32'h0000B978: begin
				q			<=			16'h0813;
		end
		32'h0000B97A: begin
				q			<=			16'h0200;
		end
		32'h0000B97C: begin
				q			<=			16'hD733;
		end
		32'h0000B97E: begin
				q			<=			16'h00E7;
		end
		32'h0000B980: begin
				q			<=			16'h0693;
		end
		32'h0000B982: begin
				q			<=			16'h0000;
		end
		32'h0000B984: begin
				q			<=			16'h8663;
		end
		32'h0000B986: begin
				q			<=			16'h0105;
		end
		32'h0000B988: begin
				q			<=			16'h0513;
		end
		32'h0000B98A: begin
				q			<=			16'h43E5;
		end
		32'h0000B98C: begin
				q			<=			16'h96B3;
		end
		32'h0000B98E: begin
				q			<=			16'h00A7;
		end
		32'h0000B990: begin
				q			<=			16'hE533;
		end
		32'h0000B992: begin
				q			<=			16'h01F6;
		end
		32'h0000B994: begin
				q			<=			16'h3533;
		end
		32'h0000B996: begin
				q			<=			16'h00A0;
		end
		32'h0000B998: begin
				q			<=			16'h6733;
		end
		32'h0000B99A: begin
				q			<=			16'h00A7;
		end
		32'h0000B99C: begin
				q			<=			16'h0793;
		end
		32'h0000B99E: begin
				q			<=			16'h0000;
		end
		32'h0000B9A0: begin
				q			<=			16'hF06F;
		end
		32'h0000B9A2: begin
				q			<=			16'hF8DF;
		end
		32'h0000B9A4: begin
				q			<=			16'h07B7;
		end
		32'h0000B9A6: begin
				q			<=			16'h0008;
		end
		32'h0000B9A8: begin
				q			<=			16'h0713;
		end
		32'h0000B9AA: begin
				q			<=			16'h0000;
		end
		32'h0000B9AC: begin
				q			<=			16'h0693;
		end
		32'h0000B9AE: begin
				q			<=			16'h7FF0;
		end
		32'h0000B9B0: begin
				q			<=			16'h0613;
		end
		32'h0000B9B2: begin
				q			<=			16'h0000;
		end
		32'h0000B9B4: begin
				q			<=			16'hF06F;
		end
		32'h0000B9B6: begin
				q			<=			16'hE85F;
		end
		32'h0000B9B8: begin
				q			<=			16'h0793;
		end
		32'h0000B9BA: begin
				q			<=			16'h0000;
		end
		32'h0000B9BC: begin
				q			<=			16'h0713;
		end
		32'h0000B9BE: begin
				q			<=			16'h0000;
		end
		32'h0000B9C0: begin
				q			<=			16'h0693;
		end
		32'h0000B9C2: begin
				q			<=			16'h7FF0;
		end
		32'h0000B9C4: begin
				q			<=			16'hF06F;
		end
		32'h0000B9C6: begin
				q			<=			16'hE75F;
		end
		32'h0000B9C8: begin
				q			<=			16'h0793;
		end
		32'h0000B9CA: begin
				q			<=			16'h0000;
		end
		32'h0000B9CC: begin
				q			<=			16'h0713;
		end
		32'h0000B9CE: begin
				q			<=			16'h0000;
		end
		32'h0000B9D0: begin
				q			<=			16'h0693;
		end
		32'h0000B9D2: begin
				q			<=			16'h0010;
		end
		32'h0000B9D4: begin
				q			<=			16'hF06F;
		end
		32'h0000B9D6: begin
				q			<=			16'hE65F;
		end
		32'h0000B9D8: begin
				q			<=			16'h0000;
		end
		32'h0000B9DA: begin
				q			<=			16'h0000;
		end
		32'h0000B9DC: begin
				q			<=			16'h0113;
		end
		32'h0000B9DE: begin
				q			<=			16'hFD01;
		end
		32'h0000B9E0: begin
				q			<=			16'h2023;
		end
		32'h0000B9E2: begin
				q			<=			16'h0321;
		end
		32'h0000B9E4: begin
				q			<=			16'h2A23;
		end
		32'h0000B9E6: begin
				q			<=			16'h0151;
		end
		32'h0000B9E8: begin
				q			<=			16'h0937;
		end
		32'h0000B9EA: begin
				q			<=			16'h0010;
		end
		32'h0000B9EC: begin
				q			<=			16'hDA93;
		end
		32'h0000B9EE: begin
				q			<=			16'h0145;
		end
		32'h0000B9F0: begin
				q			<=			16'h2E23;
		end
		32'h0000B9F2: begin
				q			<=			16'h0131;
		end
		32'h0000B9F4: begin
				q			<=			16'h2C23;
		end
		32'h0000B9F6: begin
				q			<=			16'h0141;
		end
		32'h0000B9F8: begin
				q			<=			16'h2823;
		end
		32'h0000B9FA: begin
				q			<=			16'h0161;
		end
		32'h0000B9FC: begin
				q			<=			16'h2623;
		end
		32'h0000B9FE: begin
				q			<=			16'h0171;
		end
		32'h0000BA00: begin
				q			<=			16'h0913;
		end
		32'h0000BA02: begin
				q			<=			16'hFFF9;
		end
		32'h0000BA04: begin
				q			<=			16'h2623;
		end
		32'h0000BA06: begin
				q			<=			16'h0211;
		end
		32'h0000BA08: begin
				q			<=			16'h2423;
		end
		32'h0000BA0A: begin
				q			<=			16'h0281;
		end
		32'h0000BA0C: begin
				q			<=			16'h2223;
		end
		32'h0000BA0E: begin
				q			<=			16'h0291;
		end
		32'h0000BA10: begin
				q			<=			16'hFA93;
		end
		32'h0000BA12: begin
				q			<=			16'h7FFA;
		end
		32'h0000BA14: begin
				q			<=			16'h0B13;
		end
		32'h0000BA16: begin
				q			<=			16'h0005;
		end
		32'h0000BA18: begin
				q			<=			16'h0B93;
		end
		32'h0000BA1A: begin
				q			<=			16'h0006;
		end
		32'h0000BA1C: begin
				q			<=			16'h8A13;
		end
		32'h0000BA1E: begin
				q			<=			16'h0006;
		end
		32'h0000BA20: begin
				q			<=			16'h7933;
		end
		32'h0000BA22: begin
				q			<=			16'h00B9;
		end
		32'h0000BA24: begin
				q			<=			16'hD993;
		end
		32'h0000BA26: begin
				q			<=			16'h01F5;
		end
		32'h0000BA28: begin
				q			<=			16'h8863;
		end
		32'h0000BA2A: begin
				q			<=			16'h0A0A;
		end
		32'h0000BA2C: begin
				q			<=			16'h0793;
		end
		32'h0000BA2E: begin
				q			<=			16'h7FF0;
		end
		32'h0000BA30: begin
				q			<=			16'h8663;
		end
		32'h0000BA32: begin
				q			<=			16'h10FA;
		end
		32'h0000BA34: begin
				q			<=			16'h0437;
		end
		32'h0000BA36: begin
				q			<=			16'h0080;
		end
		32'h0000BA38: begin
				q			<=			16'h1913;
		end
		32'h0000BA3A: begin
				q			<=			16'h0039;
		end
		32'h0000BA3C: begin
				q			<=			16'h6933;
		end
		32'h0000BA3E: begin
				q			<=			16'h0089;
		end
		32'h0000BA40: begin
				q			<=			16'h5413;
		end
		32'h0000BA42: begin
				q			<=			16'h01D5;
		end
		32'h0000BA44: begin
				q			<=			16'h6433;
		end
		32'h0000BA46: begin
				q			<=			16'h0124;
		end
		32'h0000BA48: begin
				q			<=			16'h1493;
		end
		32'h0000BA4A: begin
				q			<=			16'h0035;
		end
		32'h0000BA4C: begin
				q			<=			16'h8A93;
		end
		32'h0000BA4E: begin
				q			<=			16'hC01A;
		end
		32'h0000BA50: begin
				q			<=			16'h0B13;
		end
		32'h0000BA52: begin
				q			<=			16'h0000;
		end
		32'h0000BA54: begin
				q			<=			16'h5513;
		end
		32'h0000BA56: begin
				q			<=			16'h014A;
		end
		32'h0000BA58: begin
				q			<=			16'h0937;
		end
		32'h0000BA5A: begin
				q			<=			16'h0010;
		end
		32'h0000BA5C: begin
				q			<=			16'h0913;
		end
		32'h0000BA5E: begin
				q			<=			16'hFFF9;
		end
		32'h0000BA60: begin
				q			<=			16'h7513;
		end
		32'h0000BA62: begin
				q			<=			16'h7FF5;
		end
		32'h0000BA64: begin
				q			<=			16'h7933;
		end
		32'h0000BA66: begin
				q			<=			16'h0149;
		end
		32'h0000BA68: begin
				q			<=			16'h8713;
		end
		32'h0000BA6A: begin
				q			<=			16'h000B;
		end
		32'h0000BA6C: begin
				q			<=			16'h5A13;
		end
		32'h0000BA6E: begin
				q			<=			16'h01FA;
		end
		32'h0000BA70: begin
				q			<=			16'h0463;
		end
		32'h0000BA72: begin
				q			<=			16'h1005;
		end
		32'h0000BA74: begin
				q			<=			16'h0793;
		end
		32'h0000BA76: begin
				q			<=			16'h7FF0;
		end
		32'h0000BA78: begin
				q			<=			16'h0463;
		end
		32'h0000BA7A: begin
				q			<=			16'h16F5;
		end
		32'h0000BA7C: begin
				q			<=			16'h07B7;
		end
		32'h0000BA7E: begin
				q			<=			16'h0080;
		end
		32'h0000BA80: begin
				q			<=			16'h1913;
		end
		32'h0000BA82: begin
				q			<=			16'h0039;
		end
		32'h0000BA84: begin
				q			<=			16'h6933;
		end
		32'h0000BA86: begin
				q			<=			16'h00F9;
		end
		32'h0000BA88: begin
				q			<=			16'hD793;
		end
		32'h0000BA8A: begin
				q			<=			16'h01DB;
		end
		32'h0000BA8C: begin
				q			<=			16'hE7B3;
		end
		32'h0000BA8E: begin
				q			<=			16'h0127;
		end
		32'h0000BA90: begin
				q			<=			16'h9713;
		end
		32'h0000BA92: begin
				q			<=			16'h003B;
		end
		32'h0000BA94: begin
				q			<=			16'h0513;
		end
		32'h0000BA96: begin
				q			<=			16'hC015;
		end
		32'h0000BA98: begin
				q			<=			16'h0693;
		end
		32'h0000BA9A: begin
				q			<=			16'h0000;
		end
		32'h0000BA9C: begin
				q			<=			16'h1593;
		end
		32'h0000BA9E: begin
				q			<=			16'h002B;
		end
		32'h0000BAA0: begin
				q			<=			16'hE5B3;
		end
		32'h0000BAA2: begin
				q			<=			16'h00D5;
		end
		32'h0000BAA4: begin
				q			<=			16'h8533;
		end
		32'h0000BAA6: begin
				q			<=			16'h00AA;
		end
		32'h0000BAA8: begin
				q			<=			16'h8593;
		end
		32'h0000BAAA: begin
				q			<=			16'hFFF5;
		end
		32'h0000BAAC: begin
				q			<=			16'h0893;
		end
		32'h0000BAAE: begin
				q			<=			16'h00E0;
		end
		32'h0000BAB0: begin
				q			<=			16'hC633;
		end
		32'h0000BAB2: begin
				q			<=			16'h0149;
		end
		32'h0000BAB4: begin
				q			<=			16'h0813;
		end
		32'h0000BAB6: begin
				q			<=			16'h0015;
		end
		32'h0000BAB8: begin
				q			<=			16'hE063;
		end
		32'h0000BABA: begin
				q			<=			16'h16B8;
		end
		32'h0000BABC: begin
				q			<=			16'h4517;
		end
		32'h0000BABE: begin
				q			<=			16'h0000;
		end
		32'h0000BAC0: begin
				q			<=			16'h0513;
		end
		32'h0000BAC2: begin
				q			<=			16'hE385;
		end
		32'h0000BAC4: begin
				q			<=			16'h9593;
		end
		32'h0000BAC6: begin
				q			<=			16'h0025;
		end
		32'h0000BAC8: begin
				q			<=			16'h85B3;
		end
		32'h0000BACA: begin
				q			<=			16'h00A5;
		end
		32'h0000BACC: begin
				q			<=			16'hA583;
		end
		32'h0000BACE: begin
				q			<=			16'h0005;
		end
		32'h0000BAD0: begin
				q			<=			16'h85B3;
		end
		32'h0000BAD2: begin
				q			<=			16'h00A5;
		end
		32'h0000BAD4: begin
				q			<=			16'h8067;
		end
		32'h0000BAD6: begin
				q			<=			16'h0005;
		end
		32'h0000BAD8: begin
				q			<=			16'h6433;
		end
		32'h0000BADA: begin
				q			<=			16'h00A9;
		end
		32'h0000BADC: begin
				q			<=			16'h0E63;
		end
		32'h0000BADE: begin
				q			<=			16'h0604;
		end
		32'h0000BAE0: begin
				q			<=			16'h0063;
		end
		32'h0000BAE2: begin
				q			<=			16'h0409;
		end
		32'h0000BAE4: begin
				q			<=			16'h0513;
		end
		32'h0000BAE6: begin
				q			<=			16'h0009;
		end
		32'h0000BAE8: begin
				q			<=			16'h30EF;
		end
		32'h0000BAEA: begin
				q			<=			16'h5E40;
		end
		32'h0000BAEC: begin
				q			<=			16'h0793;
		end
		32'h0000BAEE: begin
				q			<=			16'hFF55;
		end
		32'h0000BAF0: begin
				q			<=			16'h0713;
		end
		32'h0000BAF2: begin
				q			<=			16'h01C0;
		end
		32'h0000BAF4: begin
				q			<=			16'h4C63;
		end
		32'h0000BAF6: begin
				q			<=			16'h02F7;
		end
		32'h0000BAF8: begin
				q			<=			16'h0413;
		end
		32'h0000BAFA: begin
				q			<=			16'h01D0;
		end
		32'h0000BAFC: begin
				q			<=			16'h0493;
		end
		32'h0000BAFE: begin
				q			<=			16'hFF85;
		end
		32'h0000BB00: begin
				q			<=			16'h0433;
		end
		32'h0000BB02: begin
				q			<=			16'h40F4;
		end
		32'h0000BB04: begin
				q			<=			16'h1933;
		end
		32'h0000BB06: begin
				q			<=			16'h0099;
		end
		32'h0000BB08: begin
				q			<=			16'h5433;
		end
		32'h0000BB0A: begin
				q			<=			16'h008B;
		end
		32'h0000BB0C: begin
				q			<=			16'h6433;
		end
		32'h0000BB0E: begin
				q			<=			16'h0124;
		end
		32'h0000BB10: begin
				q			<=			16'h14B3;
		end
		32'h0000BB12: begin
				q			<=			16'h009B;
		end
		32'h0000BB14: begin
				q			<=			16'h0A93;
		end
		32'h0000BB16: begin
				q			<=			16'hC0D0;
		end
		32'h0000BB18: begin
				q			<=			16'h8AB3;
		end
		32'h0000BB1A: begin
				q			<=			16'h40AA;
		end
		32'h0000BB1C: begin
				q			<=			16'hF06F;
		end
		32'h0000BB1E: begin
				q			<=			16'hF35F;
		end
		32'h0000BB20: begin
				q			<=			16'h30EF;
		end
		32'h0000BB22: begin
				q			<=			16'h5AC0;
		end
		32'h0000BB24: begin
				q			<=			16'h0513;
		end
		32'h0000BB26: begin
				q			<=			16'h0205;
		end
		32'h0000BB28: begin
				q			<=			16'hF06F;
		end
		32'h0000BB2A: begin
				q			<=			16'hFC5F;
		end
		32'h0000BB2C: begin
				q			<=			16'h0413;
		end
		32'h0000BB2E: begin
				q			<=			16'hFD85;
		end
		32'h0000BB30: begin
				q			<=			16'h1433;
		end
		32'h0000BB32: begin
				q			<=			16'h008B;
		end
		32'h0000BB34: begin
				q			<=			16'h0493;
		end
		32'h0000BB36: begin
				q			<=			16'h0000;
		end
		32'h0000BB38: begin
				q			<=			16'hF06F;
		end
		32'h0000BB3A: begin
				q			<=			16'hFDDF;
		end
		32'h0000BB3C: begin
				q			<=			16'h6433;
		end
		32'h0000BB3E: begin
				q			<=			16'h00A9;
		end
		32'h0000BB40: begin
				q			<=			16'h0463;
		end
		32'h0000BB42: begin
				q			<=			16'h0204;
		end
		32'h0000BB44: begin
				q			<=			16'h0493;
		end
		32'h0000BB46: begin
				q			<=			16'h0005;
		end
		32'h0000BB48: begin
				q			<=			16'h0413;
		end
		32'h0000BB4A: begin
				q			<=			16'h0009;
		end
		32'h0000BB4C: begin
				q			<=			16'h0A93;
		end
		32'h0000BB4E: begin
				q			<=			16'h7FF0;
		end
		32'h0000BB50: begin
				q			<=			16'h0B13;
		end
		32'h0000BB52: begin
				q			<=			16'h0030;
		end
		32'h0000BB54: begin
				q			<=			16'hF06F;
		end
		32'h0000BB56: begin
				q			<=			16'hF01F;
		end
		32'h0000BB58: begin
				q			<=			16'h0493;
		end
		32'h0000BB5A: begin
				q			<=			16'h0000;
		end
		32'h0000BB5C: begin
				q			<=			16'h0A93;
		end
		32'h0000BB5E: begin
				q			<=			16'h0000;
		end
		32'h0000BB60: begin
				q			<=			16'h0B13;
		end
		32'h0000BB62: begin
				q			<=			16'h0010;
		end
		32'h0000BB64: begin
				q			<=			16'hF06F;
		end
		32'h0000BB66: begin
				q			<=			16'hEF1F;
		end
		32'h0000BB68: begin
				q			<=			16'h0493;
		end
		32'h0000BB6A: begin
				q			<=			16'h0000;
		end
		32'h0000BB6C: begin
				q			<=			16'h0A93;
		end
		32'h0000BB6E: begin
				q			<=			16'h7FF0;
		end
		32'h0000BB70: begin
				q			<=			16'h0B13;
		end
		32'h0000BB72: begin
				q			<=			16'h0020;
		end
		32'h0000BB74: begin
				q			<=			16'hF06F;
		end
		32'h0000BB76: begin
				q			<=			16'hEE1F;
		end
		32'h0000BB78: begin
				q			<=			16'h67B3;
		end
		32'h0000BB7A: begin
				q			<=			16'h0179;
		end
		32'h0000BB7C: begin
				q			<=			16'h8E63;
		end
		32'h0000BB7E: begin
				q			<=			16'h0607;
		end
		32'h0000BB80: begin
				q			<=			16'h0063;
		end
		32'h0000BB82: begin
				q			<=			16'h0409;
		end
		32'h0000BB84: begin
				q			<=			16'h0513;
		end
		32'h0000BB86: begin
				q			<=			16'h0009;
		end
		32'h0000BB88: begin
				q			<=			16'h30EF;
		end
		32'h0000BB8A: begin
				q			<=			16'h5440;
		end
		32'h0000BB8C: begin
				q			<=			16'h0693;
		end
		32'h0000BB8E: begin
				q			<=			16'hFF55;
		end
		32'h0000BB90: begin
				q			<=			16'h0793;
		end
		32'h0000BB92: begin
				q			<=			16'h01C0;
		end
		32'h0000BB94: begin
				q			<=			16'hCE63;
		end
		32'h0000BB96: begin
				q			<=			16'h02D7;
		end
		32'h0000BB98: begin
				q			<=			16'h0793;
		end
		32'h0000BB9A: begin
				q			<=			16'h01D0;
		end
		32'h0000BB9C: begin
				q			<=			16'h0713;
		end
		32'h0000BB9E: begin
				q			<=			16'hFF85;
		end
		32'h0000BBA0: begin
				q			<=			16'h87B3;
		end
		32'h0000BBA2: begin
				q			<=			16'h40D7;
		end
		32'h0000BBA4: begin
				q			<=			16'h1933;
		end
		32'h0000BBA6: begin
				q			<=			16'h00E9;
		end
		32'h0000BBA8: begin
				q			<=			16'hD7B3;
		end
		32'h0000BBAA: begin
				q			<=			16'h00FB;
		end
		32'h0000BBAC: begin
				q			<=			16'hE7B3;
		end
		32'h0000BBAE: begin
				q			<=			16'h0127;
		end
		32'h0000BBB0: begin
				q			<=			16'h9733;
		end
		32'h0000BBB2: begin
				q			<=			16'h00EB;
		end
		32'h0000BBB4: begin
				q			<=			16'h0693;
		end
		32'h0000BBB6: begin
				q			<=			16'hC0D0;
		end
		32'h0000BBB8: begin
				q			<=			16'h8533;
		end
		32'h0000BBBA: begin
				q			<=			16'h40A6;
		end
		32'h0000BBBC: begin
				q			<=			16'hF06F;
		end
		32'h0000BBBE: begin
				q			<=			16'hEDDF;
		end
		32'h0000BBC0: begin
				q			<=			16'h8513;
		end
		32'h0000BBC2: begin
				q			<=			16'h000B;
		end
		32'h0000BBC4: begin
				q			<=			16'h30EF;
		end
		32'h0000BBC6: begin
				q			<=			16'h5080;
		end
		32'h0000BBC8: begin
				q			<=			16'h0513;
		end
		32'h0000BBCA: begin
				q			<=			16'h0205;
		end
		32'h0000BBCC: begin
				q			<=			16'hF06F;
		end
		32'h0000BBCE: begin
				q			<=			16'hFC1F;
		end
		32'h0000BBD0: begin
				q			<=			16'h0793;
		end
		32'h0000BBD2: begin
				q			<=			16'hFD85;
		end
		32'h0000BBD4: begin
				q			<=			16'h97B3;
		end
		32'h0000BBD6: begin
				q			<=			16'h00FB;
		end
		32'h0000BBD8: begin
				q			<=			16'h0713;
		end
		32'h0000BBDA: begin
				q			<=			16'h0000;
		end
		32'h0000BBDC: begin
				q			<=			16'hF06F;
		end
		32'h0000BBDE: begin
				q			<=			16'hFD9F;
		end
		32'h0000BBE0: begin
				q			<=			16'h67B3;
		end
		32'h0000BBE2: begin
				q			<=			16'h0179;
		end
		32'h0000BBE4: begin
				q			<=			16'h8263;
		end
		32'h0000BBE6: begin
				q			<=			16'h0207;
		end
		32'h0000BBE8: begin
				q			<=			16'h0793;
		end
		32'h0000BBEA: begin
				q			<=			16'h0009;
		end
		32'h0000BBEC: begin
				q			<=			16'h0513;
		end
		32'h0000BBEE: begin
				q			<=			16'h7FF0;
		end
		32'h0000BBF0: begin
				q			<=			16'h0693;
		end
		32'h0000BBF2: begin
				q			<=			16'h0030;
		end
		32'h0000BBF4: begin
				q			<=			16'hF06F;
		end
		32'h0000BBF6: begin
				q			<=			16'hEA9F;
		end
		32'h0000BBF8: begin
				q			<=			16'h0713;
		end
		32'h0000BBFA: begin
				q			<=			16'h0000;
		end
		32'h0000BBFC: begin
				q			<=			16'h0513;
		end
		32'h0000BBFE: begin
				q			<=			16'h0000;
		end
		32'h0000BC00: begin
				q			<=			16'h0693;
		end
		32'h0000BC02: begin
				q			<=			16'h0010;
		end
		32'h0000BC04: begin
				q			<=			16'hF06F;
		end
		32'h0000BC06: begin
				q			<=			16'hE99F;
		end
		32'h0000BC08: begin
				q			<=			16'h0713;
		end
		32'h0000BC0A: begin
				q			<=			16'h0000;
		end
		32'h0000BC0C: begin
				q			<=			16'h0513;
		end
		32'h0000BC0E: begin
				q			<=			16'h7FF0;
		end
		32'h0000BC10: begin
				q			<=			16'h0693;
		end
		32'h0000BC12: begin
				q			<=			16'h0020;
		end
		32'h0000BC14: begin
				q			<=			16'hF06F;
		end
		32'h0000BC16: begin
				q			<=			16'hE89F;
		end
		32'h0000BC18: begin
				q			<=			16'h0FB7;
		end
		32'h0000BC1A: begin
				q			<=			16'h0001;
		end
		32'h0000BC1C: begin
				q			<=			16'h8F13;
		end
		32'h0000BC1E: begin
				q			<=			16'hFFFF;
		end
		32'h0000BC20: begin
				q			<=			16'hD693;
		end
		32'h0000BC22: begin
				q			<=			16'h0104;
		end
		32'h0000BC24: begin
				q			<=			16'h5313;
		end
		32'h0000BC26: begin
				q			<=			16'h0107;
		end
		32'h0000BC28: begin
				q			<=			16'hF4B3;
		end
		32'h0000BC2A: begin
				q			<=			16'h01E4;
		end
		32'h0000BC2C: begin
				q			<=			16'h7733;
		end
		32'h0000BC2E: begin
				q			<=			16'h01E7;
		end
		32'h0000BC30: begin
				q			<=			16'h08B3;
		end
		32'h0000BC32: begin
				q			<=			16'h0293;
		end
		32'h0000BC34: begin
				q			<=			16'h85B3;
		end
		32'h0000BC36: begin
				q			<=			16'h02E4;
		end
		32'h0000BC38: begin
				q			<=			16'h82B3;
		end
		32'h0000BC3A: begin
				q			<=			16'h02E6;
		end
		32'h0000BC3C: begin
				q			<=			16'h8E33;
		end
		32'h0000BC3E: begin
				q			<=			16'h0058;
		end
		32'h0000BC40: begin
				q			<=			16'hD893;
		end
		32'h0000BC42: begin
				q			<=			16'h0105;
		end
		32'h0000BC44: begin
				q			<=			16'h88B3;
		end
		32'h0000BC46: begin
				q			<=			16'h01C8;
		end
		32'h0000BC48: begin
				q			<=			16'h8EB3;
		end
		32'h0000BC4A: begin
				q			<=			16'h0266;
		end
		32'h0000BC4C: begin
				q			<=			16'hF463;
		end
		32'h0000BC4E: begin
				q			<=			16'h0058;
		end
		32'h0000BC50: begin
				q			<=			16'h8EB3;
		end
		32'h0000BC52: begin
				q			<=			16'h01FE;
		end
		32'h0000BC54: begin
				q			<=			16'hD913;
		end
		32'h0000BC56: begin
				q			<=			16'h0108;
		end
		32'h0000BC58: begin
				q			<=			16'hF8B3;
		end
		32'h0000BC5A: begin
				q			<=			16'h01E8;
		end
		32'h0000BC5C: begin
				q			<=			16'hDF93;
		end
		32'h0000BC5E: begin
				q			<=			16'h0107;
		end
		32'h0000BC60: begin
				q			<=			16'hF5B3;
		end
		32'h0000BC62: begin
				q			<=			16'h01E5;
		end
		32'h0000BC64: begin
				q			<=			16'hF3B3;
		end
		32'h0000BC66: begin
				q			<=			16'h01E7;
		end
		32'h0000BC68: begin
				q			<=			16'h9893;
		end
		32'h0000BC6A: begin
				q			<=			16'h0108;
		end
		32'h0000BC6C: begin
				q			<=			16'h88B3;
		end
		32'h0000BC6E: begin
				q			<=			16'h00B8;
		end
		32'h0000BC70: begin
				q			<=			16'h87B3;
		end
		32'h0000BC72: begin
				q			<=			16'h0276;
		end
		32'h0000BC74: begin
				q			<=			16'h85B3;
		end
		32'h0000BC76: begin
				q			<=			16'h0293;
		end
		32'h0000BC78: begin
				q			<=			16'h84B3;
		end
		32'h0000BC7A: begin
				q			<=			16'h029F;
		end
		32'h0000BC7C: begin
				q			<=			16'h8E33;
		end
		32'h0000BC7E: begin
				q			<=			16'h00F4;
		end
		32'h0000BC80: begin
				q			<=			16'hD493;
		end
		32'h0000BC82: begin
				q			<=			16'h0105;
		end
		32'h0000BC84: begin
				q			<=			16'h84B3;
		end
		32'h0000BC86: begin
				q			<=			16'h01C4;
		end
		32'h0000BC88: begin
				q			<=			16'h86B3;
		end
		32'h0000BC8A: begin
				q			<=			16'h03F6;
		end
		32'h0000BC8C: begin
				q			<=			16'hF663;
		end
		32'h0000BC8E: begin
				q			<=			16'h00F4;
		end
		32'h0000BC90: begin
				q			<=			16'h07B7;
		end
		32'h0000BC92: begin
				q			<=			16'h0001;
		end
		32'h0000BC94: begin
				q			<=			16'h86B3;
		end
		32'h0000BC96: begin
				q			<=			16'h00F6;
		end
		32'h0000BC98: begin
				q			<=			16'hDF13;
		end
		32'h0000BC9A: begin
				q			<=			16'h0104;
		end
		32'h0000BC9C: begin
				q			<=			16'h09B7;
		end
		32'h0000BC9E: begin
				q			<=			16'h0001;
		end
		32'h0000BCA0: begin
				q			<=			16'h0F33;
		end
		32'h0000BCA2: begin
				q			<=			16'h00DF;
		end
		32'h0000BCA4: begin
				q			<=			16'h8693;
		end
		32'h0000BCA6: begin
				q			<=			16'hFFF9;
		end
		32'h0000BCA8: begin
				q			<=			16'hF4B3;
		end
		32'h0000BCAA: begin
				q			<=			16'h00D4;
		end
		32'h0000BCAC: begin
				q			<=			16'hF5B3;
		end
		32'h0000BCAE: begin
				q			<=			16'h00D5;
		end
		32'h0000BCB0: begin
				q			<=			16'h5793;
		end
		32'h0000BCB2: begin
				q			<=			16'h0104;
		end
		32'h0000BCB4: begin
				q			<=			16'h9493;
		end
		32'h0000BCB6: begin
				q			<=			16'h0104;
		end
		32'h0000BCB8: begin
				q			<=			16'h7433;
		end
		32'h0000BCBA: begin
				q			<=			16'h00D4;
		end
		32'h0000BCBC: begin
				q			<=			16'h84B3;
		end
		32'h0000BCBE: begin
				q			<=			16'h00B4;
		end
		32'h0000BCC0: begin
				q			<=			16'h06B3;
		end
		32'h0000BCC2: begin
				q			<=			16'h02E4;
		end
		32'h0000BCC4: begin
				q			<=			16'h0933;
		end
		32'h0000BCC6: begin
				q			<=			16'h0099;
		end
		32'h0000BCC8: begin
				q			<=			16'h8E33;
		end
		32'h0000BCCA: begin
				q			<=			16'h02E7;
		end
		32'h0000BCCC: begin
				q			<=			16'h05B3;
		end
		32'h0000BCCE: begin
				q			<=			16'h0283;
		end
		32'h0000BCD0: begin
				q			<=			16'h0733;
		end
		32'h0000BCD2: begin
				q			<=			16'h02F3;
		end
		32'h0000BCD4: begin
				q			<=			16'h8333;
		end
		32'h0000BCD6: begin
				q			<=			16'h01C5;
		end
		32'h0000BCD8: begin
				q			<=			16'hD593;
		end
		32'h0000BCDA: begin
				q			<=			16'h0106;
		end
		32'h0000BCDC: begin
				q			<=			16'h85B3;
		end
		32'h0000BCDE: begin
				q			<=			16'h0065;
		end
		32'h0000BCE0: begin
				q			<=			16'hF463;
		end
		32'h0000BCE2: begin
				q			<=			16'h01C5;
		end
		32'h0000BCE4: begin
				q			<=			16'h0733;
		end
		32'h0000BCE6: begin
				q			<=			16'h0137;
		end
		32'h0000BCE8: begin
				q			<=			16'hD313;
		end
		32'h0000BCEA: begin
				q			<=			16'h0105;
		end
		32'h0000BCEC: begin
				q			<=			16'h09B7;
		end
		32'h0000BCEE: begin
				q			<=			16'h0001;
		end
		32'h0000BCF0: begin
				q			<=			16'h02B3;
		end
		32'h0000BCF2: begin
				q			<=			16'h00E3;
		end
		32'h0000BCF4: begin
				q			<=			16'h8713;
		end
		32'h0000BCF6: begin
				q			<=			16'hFFF9;
		end
		32'h0000BCF8: begin
				q			<=			16'hF5B3;
		end
		32'h0000BCFA: begin
				q			<=			16'h00E5;
		end
		32'h0000BCFC: begin
				q			<=			16'hF6B3;
		end
		32'h0000BCFE: begin
				q			<=			16'h00E6;
		end
		32'h0000BD00: begin
				q			<=			16'h0333;
		end
		32'h0000BD02: begin
				q			<=			16'h0274;
		end
		32'h0000BD04: begin
				q			<=			16'h9593;
		end
		32'h0000BD06: begin
				q			<=			16'h0105;
		end
		32'h0000BD08: begin
				q			<=			16'h85B3;
		end
		32'h0000BD0A: begin
				q			<=			16'h00D5;
		end
		32'h0000BD0C: begin
				q			<=			16'h8733;
		end
		32'h0000BD0E: begin
				q			<=			16'h0277;
		end
		32'h0000BD10: begin
				q			<=			16'h8433;
		end
		32'h0000BD12: begin
				q			<=			16'h028F;
		end
		32'h0000BD14: begin
				q			<=			16'h8E33;
		end
		32'h0000BD16: begin
				q			<=			16'h02FF;
		end
		32'h0000BD18: begin
				q			<=			16'h0433;
		end
		32'h0000BD1A: begin
				q			<=			16'h00E4;
		end
		32'h0000BD1C: begin
				q			<=			16'h5793;
		end
		32'h0000BD1E: begin
				q			<=			16'h0103;
		end
		32'h0000BD20: begin
				q			<=			16'h8433;
		end
		32'h0000BD22: begin
				q			<=			16'h0087;
		end
		32'h0000BD24: begin
				q			<=			16'h7463;
		end
		32'h0000BD26: begin
				q			<=			16'h00E4;
		end
		32'h0000BD28: begin
				q			<=			16'h0E33;
		end
		32'h0000BD2A: begin
				q			<=			16'h013E;
		end
		32'h0000BD2C: begin
				q			<=			16'h07B7;
		end
		32'h0000BD2E: begin
				q			<=			16'h0001;
		end
		32'h0000BD30: begin
				q			<=			16'h8793;
		end
		32'h0000BD32: begin
				q			<=			16'hFFF7;
		end
		32'h0000BD34: begin
				q			<=			16'h76B3;
		end
		32'h0000BD36: begin
				q			<=			16'h00F4;
		end
		32'h0000BD38: begin
				q			<=			16'h7333;
		end
		32'h0000BD3A: begin
				q			<=			16'h00F3;
		end
		32'h0000BD3C: begin
				q			<=			16'h9693;
		end
		32'h0000BD3E: begin
				q			<=			16'h0106;
		end
		32'h0000BD40: begin
				q			<=			16'h8EB3;
		end
		32'h0000BD42: begin
				q			<=			16'h012E;
		end
		32'h0000BD44: begin
				q			<=			16'h86B3;
		end
		32'h0000BD46: begin
				q			<=			16'h0066;
		end
		32'h0000BD48: begin
				q			<=			16'hB4B3;
		end
		32'h0000BD4A: begin
				q			<=			16'h009E;
		end
		32'h0000BD4C: begin
				q			<=			16'h86B3;
		end
		32'h0000BD4E: begin
				q			<=			16'h01E6;
		end
		32'h0000BD50: begin
				q			<=			16'h87B3;
		end
		32'h0000BD52: begin
				q			<=			16'h0096;
		end
		32'h0000BD54: begin
				q			<=			16'h8EB3;
		end
		32'h0000BD56: begin
				q			<=			16'h00BE;
		end
		32'h0000BD58: begin
				q			<=			16'hB5B3;
		end
		32'h0000BD5A: begin
				q			<=			16'h00BE;
		end
		32'h0000BD5C: begin
				q			<=			16'h8333;
		end
		32'h0000BD5E: begin
				q			<=			16'h0057;
		end
		32'h0000BD60: begin
				q			<=			16'h0FB3;
		end
		32'h0000BD62: begin
				q			<=			16'h00B3;
		end
		32'h0000BD64: begin
				q			<=			16'hB6B3;
		end
		32'h0000BD66: begin
				q			<=			16'h01E6;
		end
		32'h0000BD68: begin
				q			<=			16'hB7B3;
		end
		32'h0000BD6A: begin
				q			<=			16'h0097;
		end
		32'h0000BD6C: begin
				q			<=			16'hE7B3;
		end
		32'h0000BD6E: begin
				q			<=			16'h00F6;
		end
		32'h0000BD70: begin
				q			<=			16'h5413;
		end
		32'h0000BD72: begin
				q			<=			16'h0104;
		end
		32'h0000BD74: begin
				q			<=			16'h3333;
		end
		32'h0000BD76: begin
				q			<=			16'h0053;
		end
		32'h0000BD78: begin
				q			<=			16'hB5B3;
		end
		32'h0000BD7A: begin
				q			<=			16'h00BF;
		end
		32'h0000BD7C: begin
				q			<=			16'h87B3;
		end
		32'h0000BD7E: begin
				q			<=			16'h0087;
		end
		32'h0000BD80: begin
				q			<=			16'h65B3;
		end
		32'h0000BD82: begin
				q			<=			16'h00B3;
		end
		32'h0000BD84: begin
				q			<=			16'h87B3;
		end
		32'h0000BD86: begin
				q			<=			16'h00B7;
		end
		32'h0000BD88: begin
				q			<=			16'h87B3;
		end
		32'h0000BD8A: begin
				q			<=			16'h01C7;
		end
		32'h0000BD8C: begin
				q			<=			16'hD713;
		end
		32'h0000BD8E: begin
				q			<=			16'h017F;
		end
		32'h0000BD90: begin
				q			<=			16'h9793;
		end
		32'h0000BD92: begin
				q			<=			16'h0097;
		end
		32'h0000BD94: begin
				q			<=			16'hE7B3;
		end
		32'h0000BD96: begin
				q			<=			16'h00E7;
		end
		32'h0000BD98: begin
				q			<=			16'h9713;
		end
		32'h0000BD9A: begin
				q			<=			16'h009E;
		end
		32'h0000BD9C: begin
				q			<=			16'h6733;
		end
		32'h0000BD9E: begin
				q			<=			16'h0117;
		end
		32'h0000BDA0: begin
				q			<=			16'h3733;
		end
		32'h0000BDA2: begin
				q			<=			16'h00E0;
		end
		32'h0000BDA4: begin
				q			<=			16'hDE93;
		end
		32'h0000BDA6: begin
				q			<=			16'h017E;
		end
		32'h0000BDA8: begin
				q			<=			16'h9693;
		end
		32'h0000BDAA: begin
				q			<=			16'h009F;
		end
		32'h0000BDAC: begin
				q			<=			16'h6733;
		end
		32'h0000BDAE: begin
				q			<=			16'h01D7;
		end
		32'h0000BDB0: begin
				q			<=			16'h6733;
		end
		32'h0000BDB2: begin
				q			<=			16'h00D7;
		end
		32'h0000BDB4: begin
				q			<=			16'h9693;
		end
		32'h0000BDB6: begin
				q			<=			16'h0077;
		end
		32'h0000BDB8: begin
				q			<=			16'hDA63;
		end
		32'h0000BDBA: begin
				q			<=			16'h1006;
		end
		32'h0000BDBC: begin
				q			<=			16'h5693;
		end
		32'h0000BDBE: begin
				q			<=			16'h0017;
		end
		32'h0000BDC0: begin
				q			<=			16'h7713;
		end
		32'h0000BDC2: begin
				q			<=			16'h0017;
		end
		32'h0000BDC4: begin
				q			<=			16'hE733;
		end
		32'h0000BDC6: begin
				q			<=			16'h00E6;
		end
		32'h0000BDC8: begin
				q			<=			16'h9693;
		end
		32'h0000BDCA: begin
				q			<=			16'h01F7;
		end
		32'h0000BDCC: begin
				q			<=			16'h6733;
		end
		32'h0000BDCE: begin
				q			<=			16'h00D7;
		end
		32'h0000BDD0: begin
				q			<=			16'hD793;
		end
		32'h0000BDD2: begin
				q			<=			16'h0017;
		end
		32'h0000BDD4: begin
				q			<=			16'h0593;
		end
		32'h0000BDD6: begin
				q			<=			16'h3FF8;
		end
		32'h0000BDD8: begin
				q			<=			16'h5E63;
		end
		32'h0000BDDA: begin
				q			<=			16'h0EB0;
		end
		32'h0000BDDC: begin
				q			<=			16'h7693;
		end
		32'h0000BDDE: begin
				q			<=			16'h0077;
		end
		32'h0000BDE0: begin
				q			<=			16'h8063;
		end
		32'h0000BDE2: begin
				q			<=			16'h0206;
		end
		32'h0000BDE4: begin
				q			<=			16'h7693;
		end
		32'h0000BDE6: begin
				q			<=			16'h00F7;
		end
		32'h0000BDE8: begin
				q			<=			16'h0513;
		end
		32'h0000BDEA: begin
				q			<=			16'h0040;
		end
		32'h0000BDEC: begin
				q			<=			16'h8A63;
		end
		32'h0000BDEE: begin
				q			<=			16'h00A6;
		end
		32'h0000BDF0: begin
				q			<=			16'h0693;
		end
		32'h0000BDF2: begin
				q			<=			16'h0047;
		end
		32'h0000BDF4: begin
				q			<=			16'hB733;
		end
		32'h0000BDF6: begin
				q			<=			16'h00E6;
		end
		32'h0000BDF8: begin
				q			<=			16'h87B3;
		end
		32'h0000BDFA: begin
				q			<=			16'h00E7;
		end
		32'h0000BDFC: begin
				q			<=			16'h8713;
		end
		32'h0000BDFE: begin
				q			<=			16'h0006;
		end
		32'h0000BE00: begin
				q			<=			16'h9693;
		end
		32'h0000BE02: begin
				q			<=			16'h0077;
		end
		32'h0000BE04: begin
				q			<=			16'hDA63;
		end
		32'h0000BE06: begin
				q			<=			16'h0006;
		end
		32'h0000BE08: begin
				q			<=			16'h06B7;
		end
		32'h0000BE0A: begin
				q			<=			16'hFF00;
		end
		32'h0000BE0C: begin
				q			<=			16'h8693;
		end
		32'h0000BE0E: begin
				q			<=			16'hFFF6;
		end
		32'h0000BE10: begin
				q			<=			16'hF7B3;
		end
		32'h0000BE12: begin
				q			<=			16'h00D7;
		end
		32'h0000BE14: begin
				q			<=			16'h0593;
		end
		32'h0000BE16: begin
				q			<=			16'h4008;
		end
		32'h0000BE18: begin
				q			<=			16'h0693;
		end
		32'h0000BE1A: begin
				q			<=			16'h7FE0;
		end
		32'h0000BE1C: begin
				q			<=			16'hCE63;
		end
		32'h0000BE1E: begin
				q			<=			16'h16B6;
		end
		32'h0000BE20: begin
				q			<=			16'h5693;
		end
		32'h0000BE22: begin
				q			<=			16'h0037;
		end
		32'h0000BE24: begin
				q			<=			16'h9713;
		end
		32'h0000BE26: begin
				q			<=			16'h01D7;
		end
		32'h0000BE28: begin
				q			<=			16'h6733;
		end
		32'h0000BE2A: begin
				q			<=			16'h00D7;
		end
		32'h0000BE2C: begin
				q			<=			16'hD793;
		end
		32'h0000BE2E: begin
				q			<=			16'h0037;
		end
		32'h0000BE30: begin
				q			<=			16'h06B7;
		end
		32'h0000BE32: begin
				q			<=			16'h0010;
		end
		32'h0000BE34: begin
				q			<=			16'h8693;
		end
		32'h0000BE36: begin
				q			<=			16'hFFF6;
		end
		32'h0000BE38: begin
				q			<=			16'hF7B3;
		end
		32'h0000BE3A: begin
				q			<=			16'h00D7;
		end
		32'h0000BE3C: begin
				q			<=			16'hF693;
		end
		32'h0000BE3E: begin
				q			<=			16'h7FF5;
		end
		32'h0000BE40: begin
				q			<=			16'h05B7;
		end
		32'h0000BE42: begin
				q			<=			16'h8010;
		end
		32'h0000BE44: begin
				q			<=			16'h8593;
		end
		32'h0000BE46: begin
				q			<=			16'hFFF5;
		end
		32'h0000BE48: begin
				q			<=			16'h9693;
		end
		32'h0000BE4A: begin
				q			<=			16'h0146;
		end
		32'h0000BE4C: begin
				q			<=			16'hF7B3;
		end
		32'h0000BE4E: begin
				q			<=			16'h00B7;
		end
		32'h0000BE50: begin
				q			<=			16'h2083;
		end
		32'h0000BE52: begin
				q			<=			16'h02C1;
		end
		32'h0000BE54: begin
				q			<=			16'h2403;
		end
		32'h0000BE56: begin
				q			<=			16'h0281;
		end
		32'h0000BE58: begin
				q			<=			16'h1613;
		end
		32'h0000BE5A: begin
				q			<=			16'h01F6;
		end
		32'h0000BE5C: begin
				q			<=			16'hE7B3;
		end
		32'h0000BE5E: begin
				q			<=			16'h00D7;
		end
		32'h0000BE60: begin
				q			<=			16'hE6B3;
		end
		32'h0000BE62: begin
				q			<=			16'h00C7;
		end
		32'h0000BE64: begin
				q			<=			16'h2483;
		end
		32'h0000BE66: begin
				q			<=			16'h0241;
		end
		32'h0000BE68: begin
				q			<=			16'h2903;
		end
		32'h0000BE6A: begin
				q			<=			16'h0201;
		end
		32'h0000BE6C: begin
				q			<=			16'h2983;
		end
		32'h0000BE6E: begin
				q			<=			16'h01C1;
		end
		32'h0000BE70: begin
				q			<=			16'h2A03;
		end
		32'h0000BE72: begin
				q			<=			16'h0181;
		end
		32'h0000BE74: begin
				q			<=			16'h2A83;
		end
		32'h0000BE76: begin
				q			<=			16'h0141;
		end
		32'h0000BE78: begin
				q			<=			16'h2B03;
		end
		32'h0000BE7A: begin
				q			<=			16'h0101;
		end
		32'h0000BE7C: begin
				q			<=			16'h2B83;
		end
		32'h0000BE7E: begin
				q			<=			16'h00C1;
		end
		32'h0000BE80: begin
				q			<=			16'h0513;
		end
		32'h0000BE82: begin
				q			<=			16'h0007;
		end
		32'h0000BE84: begin
				q			<=			16'h8593;
		end
		32'h0000BE86: begin
				q			<=			16'h0006;
		end
		32'h0000BE88: begin
				q			<=			16'h0113;
		end
		32'h0000BE8A: begin
				q			<=			16'h0301;
		end
		32'h0000BE8C: begin
				q			<=			16'h8067;
		end
		32'h0000BE8E: begin
				q			<=			16'h0000;
		end
		32'h0000BE90: begin
				q			<=			16'h8613;
		end
		32'h0000BE92: begin
				q			<=			16'h0009;
		end
		32'h0000BE94: begin
				q			<=			16'h0793;
		end
		32'h0000BE96: begin
				q			<=			16'h0004;
		end
		32'h0000BE98: begin
				q			<=			16'h8713;
		end
		32'h0000BE9A: begin
				q			<=			16'h0004;
		end
		32'h0000BE9C: begin
				q			<=			16'h0693;
		end
		32'h0000BE9E: begin
				q			<=			16'h000B;
		end
		32'h0000BEA0: begin
				q			<=			16'h0593;
		end
		32'h0000BEA2: begin
				q			<=			16'h0020;
		end
		32'h0000BEA4: begin
				q			<=			16'h8A63;
		end
		32'h0000BEA6: begin
				q			<=			16'h0EB6;
		end
		32'h0000BEA8: begin
				q			<=			16'h0593;
		end
		32'h0000BEAA: begin
				q			<=			16'h0030;
		end
		32'h0000BEAC: begin
				q			<=			16'h8C63;
		end
		32'h0000BEAE: begin
				q			<=			16'h0CB6;
		end
		32'h0000BEB0: begin
				q			<=			16'h0593;
		end
		32'h0000BEB2: begin
				q			<=			16'h0010;
		end
		32'h0000BEB4: begin
				q			<=			16'h90E3;
		end
		32'h0000BEB6: begin
				q			<=			16'hF2B6;
		end
		32'h0000BEB8: begin
				q			<=			16'h0793;
		end
		32'h0000BEBA: begin
				q			<=			16'h0000;
		end
		32'h0000BEBC: begin
				q			<=			16'h0713;
		end
		32'h0000BEBE: begin
				q			<=			16'h0000;
		end
		32'h0000BEC0: begin
				q			<=			16'h006F;
		end
		32'h0000BEC2: begin
				q			<=			16'h0880;
		end
		32'h0000BEC4: begin
				q			<=			16'h0613;
		end
		32'h0000BEC6: begin
				q			<=			16'h000A;
		end
		32'h0000BEC8: begin
				q			<=			16'hF06F;
		end
		32'h0000BECA: begin
				q			<=			16'hFD9F;
		end
		32'h0000BECC: begin
				q			<=			16'h0813;
		end
		32'h0000BECE: begin
				q			<=			16'h0005;
		end
		32'h0000BED0: begin
				q			<=			16'hF06F;
		end
		32'h0000BED2: begin
				q			<=			16'hF05F;
		end
		32'h0000BED4: begin
				q			<=			16'h0513;
		end
		32'h0000BED6: begin
				q			<=			16'h0010;
		end
		32'h0000BED8: begin
				q			<=			16'h0533;
		end
		32'h0000BEDA: begin
				q			<=			16'h40B5;
		end
		32'h0000BEDC: begin
				q			<=			16'h0693;
		end
		32'h0000BEDE: begin
				q			<=			16'h0380;
		end
		32'h0000BEE0: begin
				q			<=			16'hCCE3;
		end
		32'h0000BEE2: begin
				q			<=			16'hFCA6;
		end
		32'h0000BEE4: begin
				q			<=			16'h0693;
		end
		32'h0000BEE6: begin
				q			<=			16'h01F0;
		end
		32'h0000BEE8: begin
				q			<=			16'hC463;
		end
		32'h0000BEEA: begin
				q			<=			16'h06A6;
		end
		32'h0000BEEC: begin
				q			<=			16'h0813;
		end
		32'h0000BEEE: begin
				q			<=			16'h41E8;
		end
		32'h0000BEF0: begin
				q			<=			16'h96B3;
		end
		32'h0000BEF2: begin
				q			<=			16'h0107;
		end
		32'h0000BEF4: begin
				q			<=			16'h55B3;
		end
		32'h0000BEF6: begin
				q			<=			16'h00A7;
		end
		32'h0000BEF8: begin
				q			<=			16'h1733;
		end
		32'h0000BEFA: begin
				q			<=			16'h0107;
		end
		32'h0000BEFC: begin
				q			<=			16'hE6B3;
		end
		32'h0000BEFE: begin
				q			<=			16'h00B6;
		end
		32'h0000BF00: begin
				q			<=			16'h3733;
		end
		32'h0000BF02: begin
				q			<=			16'h00E0;
		end
		32'h0000BF04: begin
				q			<=			16'hE733;
		end
		32'h0000BF06: begin
				q			<=			16'h00E6;
		end
		32'h0000BF08: begin
				q			<=			16'hD7B3;
		end
		32'h0000BF0A: begin
				q			<=			16'h00A7;
		end
		32'h0000BF0C: begin
				q			<=			16'h7693;
		end
		32'h0000BF0E: begin
				q			<=			16'h0077;
		end
		32'h0000BF10: begin
				q			<=			16'h8063;
		end
		32'h0000BF12: begin
				q			<=			16'h0206;
		end
		32'h0000BF14: begin
				q			<=			16'h7693;
		end
		32'h0000BF16: begin
				q			<=			16'h00F7;
		end
		32'h0000BF18: begin
				q			<=			16'h0593;
		end
		32'h0000BF1A: begin
				q			<=			16'h0040;
		end
		32'h0000BF1C: begin
				q			<=			16'h8A63;
		end
		32'h0000BF1E: begin
				q			<=			16'h00B6;
		end
		32'h0000BF20: begin
				q			<=			16'h0693;
		end
		32'h0000BF22: begin
				q			<=			16'h0047;
		end
		32'h0000BF24: begin
				q			<=			16'hB733;
		end
		32'h0000BF26: begin
				q			<=			16'h00E6;
		end
		32'h0000BF28: begin
				q			<=			16'h87B3;
		end
		32'h0000BF2A: begin
				q			<=			16'h00E7;
		end
		32'h0000BF2C: begin
				q			<=			16'h8713;
		end
		32'h0000BF2E: begin
				q			<=			16'h0006;
		end
		32'h0000BF30: begin
				q			<=			16'h9693;
		end
		32'h0000BF32: begin
				q			<=			16'h0087;
		end
		32'h0000BF34: begin
				q			<=			16'hCA63;
		end
		32'h0000BF36: begin
				q			<=			16'h0606;
		end
		32'h0000BF38: begin
				q			<=			16'h9693;
		end
		32'h0000BF3A: begin
				q			<=			16'h01D7;
		end
		32'h0000BF3C: begin
				q			<=			16'h5713;
		end
		32'h0000BF3E: begin
				q			<=			16'h0037;
		end
		32'h0000BF40: begin
				q			<=			16'hE733;
		end
		32'h0000BF42: begin
				q			<=			16'h00E6;
		end
		32'h0000BF44: begin
				q			<=			16'hD793;
		end
		32'h0000BF46: begin
				q			<=			16'h0037;
		end
		32'h0000BF48: begin
				q			<=			16'h0593;
		end
		32'h0000BF4A: begin
				q			<=			16'h0000;
		end
		32'h0000BF4C: begin
				q			<=			16'hF06F;
		end
		32'h0000BF4E: begin
				q			<=			16'hEE5F;
		end
		32'h0000BF50: begin
				q			<=			16'h0693;
		end
		32'h0000BF52: begin
				q			<=			16'hFE10;
		end
		32'h0000BF54: begin
				q			<=			16'h86B3;
		end
		32'h0000BF56: begin
				q			<=			16'h40B6;
		end
		32'h0000BF58: begin
				q			<=			16'h0893;
		end
		32'h0000BF5A: begin
				q			<=			16'h0200;
		end
		32'h0000BF5C: begin
				q			<=			16'hD6B3;
		end
		32'h0000BF5E: begin
				q			<=			16'h00D7;
		end
		32'h0000BF60: begin
				q			<=			16'h0593;
		end
		32'h0000BF62: begin
				q			<=			16'h0000;
		end
		32'h0000BF64: begin
				q			<=			16'h0663;
		end
		32'h0000BF66: begin
				q			<=			16'h0115;
		end
		32'h0000BF68: begin
				q			<=			16'h0813;
		end
		32'h0000BF6A: begin
				q			<=			16'h43E8;
		end
		32'h0000BF6C: begin
				q			<=			16'h95B3;
		end
		32'h0000BF6E: begin
				q			<=			16'h0107;
		end
		32'h0000BF70: begin
				q			<=			16'hE733;
		end
		32'h0000BF72: begin
				q			<=			16'h00E5;
		end
		32'h0000BF74: begin
				q			<=			16'h3733;
		end
		32'h0000BF76: begin
				q			<=			16'h00E0;
		end
		32'h0000BF78: begin
				q			<=			16'hE733;
		end
		32'h0000BF7A: begin
				q			<=			16'h00E6;
		end
		32'h0000BF7C: begin
				q			<=			16'h0793;
		end
		32'h0000BF7E: begin
				q			<=			16'h0000;
		end
		32'h0000BF80: begin
				q			<=			16'hF06F;
		end
		32'h0000BF82: begin
				q			<=			16'hF8DF;
		end
		32'h0000BF84: begin
				q			<=			16'h07B7;
		end
		32'h0000BF86: begin
				q			<=			16'h0008;
		end
		32'h0000BF88: begin
				q			<=			16'h0713;
		end
		32'h0000BF8A: begin
				q			<=			16'h0000;
		end
		32'h0000BF8C: begin
				q			<=			16'h0593;
		end
		32'h0000BF8E: begin
				q			<=			16'h7FF0;
		end
		32'h0000BF90: begin
				q			<=			16'h0613;
		end
		32'h0000BF92: begin
				q			<=			16'h0000;
		end
		32'h0000BF94: begin
				q			<=			16'hF06F;
		end
		32'h0000BF96: begin
				q			<=			16'hE9DF;
		end
		32'h0000BF98: begin
				q			<=			16'h0793;
		end
		32'h0000BF9A: begin
				q			<=			16'h0000;
		end
		32'h0000BF9C: begin
				q			<=			16'h0713;
		end
		32'h0000BF9E: begin
				q			<=			16'h0000;
		end
		32'h0000BFA0: begin
				q			<=			16'h0593;
		end
		32'h0000BFA2: begin
				q			<=			16'h7FF0;
		end
		32'h0000BFA4: begin
				q			<=			16'hF06F;
		end
		32'h0000BFA6: begin
				q			<=			16'hE8DF;
		end
		32'h0000BFA8: begin
				q			<=			16'h0793;
		end
		32'h0000BFAA: begin
				q			<=			16'h0000;
		end
		32'h0000BFAC: begin
				q			<=			16'h0713;
		end
		32'h0000BFAE: begin
				q			<=			16'h0000;
		end
		32'h0000BFB0: begin
				q			<=			16'h0593;
		end
		32'h0000BFB2: begin
				q			<=			16'h0010;
		end
		32'h0000BFB4: begin
				q			<=			16'hF06F;
		end
		32'h0000BFB6: begin
				q			<=			16'hE7DF;
		end
		32'h0000BFB8: begin
				q			<=			16'h0000;
		end
		32'h0000BFBA: begin
				q			<=			16'h0000;
		end
		32'h0000BFBC: begin
				q			<=			16'h2783;
		end
		32'h0000BFBE: begin
				q			<=			16'h00C5;
		end
		32'h0000BFC0: begin
				q			<=			16'hAF03;
		end
		32'h0000BFC2: begin
				q			<=			16'h0005;
		end
		32'h0000BFC4: begin
				q			<=			16'hAF83;
		end
		32'h0000BFC6: begin
				q			<=			16'h0045;
		end
		32'h0000BFC8: begin
				q			<=			16'hA283;
		end
		32'h0000BFCA: begin
				q			<=			16'h0085;
		end
		32'h0000BFCC: begin
				q			<=			16'hA583;
		end
		32'h0000BFCE: begin
				q			<=			16'h00C5;
		end
		32'h0000BFD0: begin
				q			<=			16'h8737;
		end
		32'h0000BFD2: begin
				q			<=			16'h0000;
		end
		32'h0000BFD4: begin
				q			<=			16'hD693;
		end
		32'h0000BFD6: begin
				q			<=			16'h0107;
		end
		32'h0000BFD8: begin
				q			<=			16'h0713;
		end
		32'h0000BFDA: begin
				q			<=			16'hFFF7;
		end
		32'h0000BFDC: begin
				q			<=			16'h9813;
		end
		32'h0000BFDE: begin
				q			<=			16'h0107;
		end
		32'h0000BFE0: begin
				q			<=			16'h9E93;
		end
		32'h0000BFE2: begin
				q			<=			16'h0105;
		end
		32'h0000BFE4: begin
				q			<=			16'hD613;
		end
		32'h0000BFE6: begin
				q			<=			16'h01F7;
		end
		32'h0000BFE8: begin
				q			<=			16'h76B3;
		end
		32'h0000BFEA: begin
				q			<=			16'h00D7;
		end
		32'h0000BFEC: begin
				q			<=			16'hD793;
		end
		32'h0000BFEE: begin
				q			<=			16'h0105;
		end
		32'h0000BFF0: begin
				q			<=			16'h0113;
		end
		32'h0000BFF2: begin
				q			<=			16'hFF01;
		end
		32'h0000BFF4: begin
				q			<=			16'h2883;
		end
		32'h0000BFF6: begin
				q			<=			16'h0005;
		end
		32'h0000BFF8: begin
				q			<=			16'h2303;
		end
		32'h0000BFFA: begin
				q			<=			16'h0045;
		end
		32'h0000BFFC: begin
				q			<=			16'h2E03;
		end
		32'h0000BFFE: begin
				q			<=			16'h0085;
		end
		32'h0000C000: begin
				q			<=			16'h5813;
		end
		32'h0000C002: begin
				q			<=			16'h0108;
		end
		32'h0000C004: begin
				q			<=			16'hDE93;
		end
		32'h0000C006: begin
				q			<=			16'h010E;
		end
		32'h0000C008: begin
				q			<=			16'h77B3;
		end
		32'h0000C00A: begin
				q			<=			16'h00F7;
		end
		32'h0000C00C: begin
				q			<=			16'hD593;
		end
		32'h0000C00E: begin
				q			<=			16'h01F5;
		end
		32'h0000C010: begin
				q			<=			16'h9063;
		end
		32'h0000C012: begin
				q			<=			16'h02E6;
		end
		32'h0000C014: begin
				q			<=			16'hE733;
		end
		32'h0000C016: begin
				q			<=			16'h0068;
		end
		32'h0000C018: begin
				q			<=			16'h6733;
		end
		32'h0000C01A: begin
				q			<=			16'h01C7;
		end
		32'h0000C01C: begin
				q			<=			16'h6733;
		end
		32'h0000C01E: begin
				q			<=			16'h0107;
		end
		32'h0000C020: begin
				q			<=			16'h0513;
		end
		32'h0000C022: begin
				q			<=			16'h0010;
		end
		32'h0000C024: begin
				q			<=			16'h1A63;
		end
		32'h0000C026: begin
				q			<=			16'h0407;
		end
		32'h0000C028: begin
				q			<=			16'h9863;
		end
		32'h0000C02A: begin
				q			<=			16'h04D7;
		end
		32'h0000C02C: begin
				q			<=			16'h006F;
		end
		32'h0000C02E: begin
				q			<=			16'h0080;
		end
		32'h0000C030: begin
				q			<=			16'h9C63;
		end
		32'h0000C032: begin
				q			<=			16'h00E7;
		end
		32'h0000C034: begin
				q			<=			16'h6733;
		end
		32'h0000C036: begin
				q			<=			16'h01FF;
		end
		32'h0000C038: begin
				q			<=			16'h6733;
		end
		32'h0000C03A: begin
				q			<=			16'h0057;
		end
		32'h0000C03C: begin
				q			<=			16'h6733;
		end
		32'h0000C03E: begin
				q			<=			16'h01D7;
		end
		32'h0000C040: begin
				q			<=			16'h0513;
		end
		32'h0000C042: begin
				q			<=			16'h0010;
		end
		32'h0000C044: begin
				q			<=			16'h1A63;
		end
		32'h0000C046: begin
				q			<=			16'h0207;
		end
		32'h0000C048: begin
				q			<=			16'h0513;
		end
		32'h0000C04A: begin
				q			<=			16'h0010;
		end
		32'h0000C04C: begin
				q			<=			16'h9663;
		end
		32'h0000C04E: begin
				q			<=			16'h02D7;
		end
		32'h0000C050: begin
				q			<=			16'h9463;
		end
		32'h0000C052: begin
				q			<=			16'h03E8;
		end
		32'h0000C054: begin
				q			<=			16'h1263;
		end
		32'h0000C056: begin
				q			<=			16'h03F3;
		end
		32'h0000C058: begin
				q			<=			16'h1063;
		end
		32'h0000C05A: begin
				q			<=			16'h025E;
		end
		32'h0000C05C: begin
				q			<=			16'h1E63;
		end
		32'h0000C05E: begin
				q			<=			16'h01D8;
		end
		32'h0000C060: begin
				q			<=			16'h0063;
		end
		32'h0000C062: begin
				q			<=			16'h02B6;
		end
		32'h0000C064: begin
				q			<=			16'h9A63;
		end
		32'h0000C066: begin
				q			<=			16'h0007;
		end
		32'h0000C068: begin
				q			<=			16'hE533;
		end
		32'h0000C06A: begin
				q			<=			16'h0068;
		end
		32'h0000C06C: begin
				q			<=			16'h6533;
		end
		32'h0000C06E: begin
				q			<=			16'h01C5;
		end
		32'h0000C070: begin
				q			<=			16'h6533;
		end
		32'h0000C072: begin
				q			<=			16'h0105;
		end
		32'h0000C074: begin
				q			<=			16'h3533;
		end
		32'h0000C076: begin
				q			<=			16'h00A0;
		end
		32'h0000C078: begin
				q			<=			16'h0113;
		end
		32'h0000C07A: begin
				q			<=			16'h0101;
		end
		32'h0000C07C: begin
				q			<=			16'h8067;
		end
		32'h0000C07E: begin
				q			<=			16'h0000;
		end
		32'h0000C080: begin
				q			<=			16'h0513;
		end
		32'h0000C082: begin
				q			<=			16'h0000;
		end
		32'h0000C084: begin
				q			<=			16'hF06F;
		end
		32'h0000C086: begin
				q			<=			16'hFF5F;
		end
		32'h0000C088: begin
				q			<=			16'h0000;
		end
		32'h0000C08A: begin
				q			<=			16'h0000;
		end
		32'h0000C08C: begin
				q			<=			16'h2783;
		end
		32'h0000C08E: begin
				q			<=			16'h00C5;
		end
		32'h0000C090: begin
				q			<=			16'hA883;
		end
		32'h0000C092: begin
				q			<=			16'h00C5;
		end
		32'h0000C094: begin
				q			<=			16'h2F03;
		end
		32'h0000C096: begin
				q			<=			16'h0005;
		end
		32'h0000C098: begin
				q			<=			16'h2603;
		end
		32'h0000C09A: begin
				q			<=			16'h0045;
		end
		32'h0000C09C: begin
				q			<=			16'h2803;
		end
		32'h0000C09E: begin
				q			<=			16'h0085;
		end
		32'h0000C0A0: begin
				q			<=			16'h8537;
		end
		32'h0000C0A2: begin
				q			<=			16'h0000;
		end
		32'h0000C0A4: begin
				q			<=			16'hD713;
		end
		32'h0000C0A6: begin
				q			<=			16'h0107;
		end
		32'h0000C0A8: begin
				q			<=			16'h0513;
		end
		32'h0000C0AA: begin
				q			<=			16'hFFF5;
		end
		32'h0000C0AC: begin
				q			<=			16'h9E93;
		end
		32'h0000C0AE: begin
				q			<=			16'h0108;
		end
		32'h0000C0B0: begin
				q			<=			16'hD693;
		end
		32'h0000C0B2: begin
				q			<=			16'h0108;
		end
		32'h0000C0B4: begin
				q			<=			16'hA283;
		end
		32'h0000C0B6: begin
				q			<=			16'h0005;
		end
		32'h0000C0B8: begin
				q			<=			16'hA303;
		end
		32'h0000C0BA: begin
				q			<=			16'h0045;
		end
		32'h0000C0BC: begin
				q			<=			16'hAE03;
		end
		32'h0000C0BE: begin
				q			<=			16'h0085;
		end
		32'h0000C0C0: begin
				q			<=			16'h7733;
		end
		32'h0000C0C2: begin
				q			<=			16'h00E5;
		end
		32'h0000C0C4: begin
				q			<=			16'h9593;
		end
		32'h0000C0C6: begin
				q			<=			16'h0107;
		end
		32'h0000C0C8: begin
				q			<=			16'h0113;
		end
		32'h0000C0CA: begin
				q			<=			16'hFF01;
		end
		32'h0000C0CC: begin
				q			<=			16'hD593;
		end
		32'h0000C0CE: begin
				q			<=			16'h0105;
		end
		32'h0000C0D0: begin
				q			<=			16'hD793;
		end
		32'h0000C0D2: begin
				q			<=			16'h01F7;
		end
		32'h0000C0D4: begin
				q			<=			16'hDE93;
		end
		32'h0000C0D6: begin
				q			<=			16'h010E;
		end
		32'h0000C0D8: begin
				q			<=			16'h76B3;
		end
		32'h0000C0DA: begin
				q			<=			16'h00D5;
		end
		32'h0000C0DC: begin
				q			<=			16'hD893;
		end
		32'h0000C0DE: begin
				q			<=			16'h01F8;
		end
		32'h0000C0E0: begin
				q			<=			16'h1063;
		end
		32'h0000C0E2: begin
				q			<=			16'h02A7;
		end
		32'h0000C0E4: begin
				q			<=			16'h6FB3;
		end
		32'h0000C0E6: begin
				q			<=			16'h00CF;
		end
		32'h0000C0E8: begin
				q			<=			16'hEFB3;
		end
		32'h0000C0EA: begin
				q			<=			16'h010F;
		end
		32'h0000C0EC: begin
				q			<=			16'hEFB3;
		end
		32'h0000C0EE: begin
				q			<=			16'h00BF;
		end
		32'h0000C0F0: begin
				q			<=			16'h0513;
		end
		32'h0000C0F2: begin
				q			<=			16'hFFE0;
		end
		32'h0000C0F4: begin
				q			<=			16'h8063;
		end
		32'h0000C0F6: begin
				q			<=			16'h0E0F;
		end
		32'h0000C0F8: begin
				q			<=			16'h0113;
		end
		32'h0000C0FA: begin
				q			<=			16'h0101;
		end
		32'h0000C0FC: begin
				q			<=			16'h8067;
		end
		32'h0000C0FE: begin
				q			<=			16'h0000;
		end
		32'h0000C100: begin
				q			<=			16'h9863;
		end
		32'h0000C102: begin
				q			<=			16'h02A6;
		end
		32'h0000C104: begin
				q			<=			16'hEFB3;
		end
		32'h0000C106: begin
				q			<=			16'h0062;
		end
		32'h0000C108: begin
				q			<=			16'hEFB3;
		end
		32'h0000C10A: begin
				q			<=			16'h01CF;
		end
		32'h0000C10C: begin
				q			<=			16'hEFB3;
		end
		32'h0000C10E: begin
				q			<=			16'h01DF;
		end
		32'h0000C110: begin
				q			<=			16'h0513;
		end
		32'h0000C112: begin
				q			<=			16'hFFE0;
		end
		32'h0000C114: begin
				q			<=			16'h92E3;
		end
		32'h0000C116: begin
				q			<=			16'hFE0F;
		end
		32'h0000C118: begin
				q			<=			16'h1263;
		end
		32'h0000C11A: begin
				q			<=			16'h0407;
		end
		32'h0000C11C: begin
				q			<=			16'h6533;
		end
		32'h0000C11E: begin
				q			<=			16'h00CF;
		end
		32'h0000C120: begin
				q			<=			16'h6533;
		end
		32'h0000C122: begin
				q			<=			16'h0105;
		end
		32'h0000C124: begin
				q			<=			16'h6533;
		end
		32'h0000C126: begin
				q			<=			16'h00B5;
		end
		32'h0000C128: begin
				q			<=			16'h3513;
		end
		32'h0000C12A: begin
				q			<=			16'h0015;
		end
		32'h0000C12C: begin
				q			<=			16'h006F;
		end
		32'h0000C12E: begin
				q			<=			16'h02C0;
		end
		32'h0000C130: begin
				q			<=			16'h1463;
		end
		32'h0000C132: begin
				q			<=			16'h0A07;
		end
		32'h0000C134: begin
				q			<=			16'h6533;
		end
		32'h0000C136: begin
				q			<=			16'h00CF;
		end
		32'h0000C138: begin
				q			<=			16'h6533;
		end
		32'h0000C13A: begin
				q			<=			16'h0105;
		end
		32'h0000C13C: begin
				q			<=			16'h6533;
		end
		32'h0000C13E: begin
				q			<=			16'h00B5;
		end
		32'h0000C140: begin
				q			<=			16'h3513;
		end
		32'h0000C142: begin
				q			<=			16'h0015;
		end
		32'h0000C144: begin
				q			<=			16'h9A63;
		end
		32'h0000C146: begin
				q			<=			16'h0006;
		end
		32'h0000C148: begin
				q			<=			16'hEFB3;
		end
		32'h0000C14A: begin
				q			<=			16'h0062;
		end
		32'h0000C14C: begin
				q			<=			16'hEFB3;
		end
		32'h0000C14E: begin
				q			<=			16'h01CF;
		end
		32'h0000C150: begin
				q			<=			16'hEFB3;
		end
		32'h0000C152: begin
				q			<=			16'h01DF;
		end
		32'h0000C154: begin
				q			<=			16'h8C63;
		end
		32'h0000C156: begin
				q			<=			16'h060F;
		end
		32'h0000C158: begin
				q			<=			16'h1A63;
		end
		32'h0000C15A: begin
				q			<=			16'h0005;
		end
		32'h0000C15C: begin
				q			<=			16'h8E63;
		end
		32'h0000C15E: begin
				q			<=			16'h0117;
		end
		32'h0000C160: begin
				q			<=			16'h0513;
		end
		32'h0000C162: begin
				q			<=			16'h0010;
		end
		32'h0000C164: begin
				q			<=			16'h8AE3;
		end
		32'h0000C166: begin
				q			<=			16'hF807;
		end
		32'h0000C168: begin
				q			<=			16'h006F;
		end
		32'h0000C16A: begin
				q			<=			16'h0080;
		end
		32'h0000C16C: begin
				q			<=			16'h96E3;
		end
		32'h0000C16E: begin
				q			<=			16'hF808;
		end
		32'h0000C170: begin
				q			<=			16'h0513;
		end
		32'h0000C172: begin
				q			<=			16'hFFF0;
		end
		32'h0000C174: begin
				q			<=			16'hF06F;
		end
		32'h0000C176: begin
				q			<=			16'hF85F;
		end
		32'h0000C178: begin
				q			<=			16'hC4E3;
		end
		32'h0000C17A: begin
				q			<=			16'hFEE6;
		end
		32'h0000C17C: begin
				q			<=			16'h5A63;
		end
		32'h0000C17E: begin
				q			<=			16'h00D7;
		end
		32'h0000C180: begin
				q			<=			16'h0513;
		end
		32'h0000C182: begin
				q			<=			16'hFFF0;
		end
		32'h0000C184: begin
				q			<=			16'h8AE3;
		end
		32'h0000C186: begin
				q			<=			16'hF607;
		end
		32'h0000C188: begin
				q			<=			16'h0513;
		end
		32'h0000C18A: begin
				q			<=			16'h0010;
		end
		32'h0000C18C: begin
				q			<=			16'hF06F;
		end
		32'h0000C18E: begin
				q			<=			16'hF6DF;
		end
		32'h0000C190: begin
				q			<=			16'hE8E3;
		end
		32'h0000C192: begin
				q			<=			16'hFCBE;
		end
		32'h0000C194: begin
				q			<=			16'h9663;
		end
		32'h0000C196: begin
				q			<=			16'h03D5;
		end
		32'h0000C198: begin
				q			<=			16'h64E3;
		end
		32'h0000C19A: begin
				q			<=			16'hFD0E;
		end
		32'h0000C19C: begin
				q			<=			16'h1463;
		end
		32'h0000C19E: begin
				q			<=			16'h05C8;
		end
		32'h0000C1A0: begin
				q			<=			16'h60E3;
		end
		32'h0000C1A2: begin
				q			<=			16'hFCC3;
		end
		32'h0000C1A4: begin
				q			<=			16'h1463;
		end
		32'h0000C1A6: begin
				q			<=			16'h0066;
		end
		32'h0000C1A8: begin
				q			<=			16'hECE3;
		end
		32'h0000C1AA: begin
				q			<=			16'hFBE2;
		end
		32'h0000C1AC: begin
				q			<=			16'h6AE3;
		end
		32'h0000C1AE: begin
				q			<=			16'hFC66;
		end
		32'h0000C1B0: begin
				q			<=			16'h0513;
		end
		32'h0000C1B2: begin
				q			<=			16'h0000;
		end
		32'h0000C1B4: begin
				q			<=			16'h12E3;
		end
		32'h0000C1B6: begin
				q			<=			16'hF466;
		end
		32'h0000C1B8: begin
				q			<=			16'h64E3;
		end
		32'h0000C1BA: begin
				q			<=			16'hFC5F;
		end
		32'h0000C1BC: begin
				q			<=			16'hF06F;
		end
		32'h0000C1BE: begin
				q			<=			16'hF3DF;
		end
		32'h0000C1C0: begin
				q			<=			16'hE0E3;
		end
		32'h0000C1C2: begin
				q			<=			16'hFDD5;
		end
		32'h0000C1C4: begin
				q			<=			16'h0513;
		end
		32'h0000C1C6: begin
				q			<=			16'h0000;
		end
		32'h0000C1C8: begin
				q			<=			16'hF06F;
		end
		32'h0000C1CA: begin
				q			<=			16'hF31F;
		end
		32'h0000C1CC: begin
				q			<=			16'h1CE3;
		end
		32'h0000C1CE: begin
				q			<=			16'hFE05;
		end
		32'h0000C1D0: begin
				q			<=			16'hF06F;
		end
		32'h0000C1D2: begin
				q			<=			16'hF91F;
		end
		32'h0000C1D4: begin
				q			<=			16'h88E3;
		end
		32'h0000C1D6: begin
				q			<=			16'hF2E6;
		end
		32'h0000C1D8: begin
				q			<=			16'h0513;
		end
		32'h0000C1DA: begin
				q			<=			16'h0000;
		end
		32'h0000C1DC: begin
				q			<=			16'h86E3;
		end
		32'h0000C1DE: begin
				q			<=			16'hF606;
		end
		32'h0000C1E0: begin
				q			<=			16'hF06F;
		end
		32'h0000C1E2: begin
				q			<=			16'hF7DF;
		end
		32'h0000C1E4: begin
				q			<=			16'h6EE3;
		end
		32'h0000C1E6: begin
				q			<=			16'hF9C8;
		end
		32'h0000C1E8: begin
				q			<=			16'hF06F;
		end
		32'h0000C1EA: begin
				q			<=			16'hFDDF;
		end
		32'h0000C1EC: begin
				q			<=			16'h0000;
		end
		32'h0000C1EE: begin
				q			<=			16'h0000;
		end
		32'h0000C1F0: begin
				q			<=			16'h2783;
		end
		32'h0000C1F2: begin
				q			<=			16'h00C5;
		end
		32'h0000C1F4: begin
				q			<=			16'hA883;
		end
		32'h0000C1F6: begin
				q			<=			16'h00C5;
		end
		32'h0000C1F8: begin
				q			<=			16'h2F03;
		end
		32'h0000C1FA: begin
				q			<=			16'h0005;
		end
		32'h0000C1FC: begin
				q			<=			16'h2603;
		end
		32'h0000C1FE: begin
				q			<=			16'h0045;
		end
		32'h0000C200: begin
				q			<=			16'h2803;
		end
		32'h0000C202: begin
				q			<=			16'h0085;
		end
		32'h0000C204: begin
				q			<=			16'h8537;
		end
		32'h0000C206: begin
				q			<=			16'h0000;
		end
		32'h0000C208: begin
				q			<=			16'hD713;
		end
		32'h0000C20A: begin
				q			<=			16'h0107;
		end
		32'h0000C20C: begin
				q			<=			16'h0513;
		end
		32'h0000C20E: begin
				q			<=			16'hFFF5;
		end
		32'h0000C210: begin
				q			<=			16'h9E93;
		end
		32'h0000C212: begin
				q			<=			16'h0108;
		end
		32'h0000C214: begin
				q			<=			16'hD693;
		end
		32'h0000C216: begin
				q			<=			16'h0108;
		end
		32'h0000C218: begin
				q			<=			16'hA283;
		end
		32'h0000C21A: begin
				q			<=			16'h0005;
		end
		32'h0000C21C: begin
				q			<=			16'hA303;
		end
		32'h0000C21E: begin
				q			<=			16'h0045;
		end
		32'h0000C220: begin
				q			<=			16'hAE03;
		end
		32'h0000C222: begin
				q			<=			16'h0085;
		end
		32'h0000C224: begin
				q			<=			16'h7733;
		end
		32'h0000C226: begin
				q			<=			16'h00E5;
		end
		32'h0000C228: begin
				q			<=			16'h9593;
		end
		32'h0000C22A: begin
				q			<=			16'h0107;
		end
		32'h0000C22C: begin
				q			<=			16'h0113;
		end
		32'h0000C22E: begin
				q			<=			16'hFF01;
		end
		32'h0000C230: begin
				q			<=			16'hD593;
		end
		32'h0000C232: begin
				q			<=			16'h0105;
		end
		32'h0000C234: begin
				q			<=			16'hD793;
		end
		32'h0000C236: begin
				q			<=			16'h01F7;
		end
		32'h0000C238: begin
				q			<=			16'hDE93;
		end
		32'h0000C23A: begin
				q			<=			16'h010E;
		end
		32'h0000C23C: begin
				q			<=			16'h76B3;
		end
		32'h0000C23E: begin
				q			<=			16'h00D5;
		end
		32'h0000C240: begin
				q			<=			16'hD893;
		end
		32'h0000C242: begin
				q			<=			16'h01F8;
		end
		32'h0000C244: begin
				q			<=			16'h1063;
		end
		32'h0000C246: begin
				q			<=			16'h02A7;
		end
		32'h0000C248: begin
				q			<=			16'h6FB3;
		end
		32'h0000C24A: begin
				q			<=			16'h00CF;
		end
		32'h0000C24C: begin
				q			<=			16'hEFB3;
		end
		32'h0000C24E: begin
				q			<=			16'h010F;
		end
		32'h0000C250: begin
				q			<=			16'hEFB3;
		end
		32'h0000C252: begin
				q			<=			16'h00BF;
		end
		32'h0000C254: begin
				q			<=			16'h0513;
		end
		32'h0000C256: begin
				q			<=			16'h0020;
		end
		32'h0000C258: begin
				q			<=			16'h8063;
		end
		32'h0000C25A: begin
				q			<=			16'h0E0F;
		end
		32'h0000C25C: begin
				q			<=			16'h0113;
		end
		32'h0000C25E: begin
				q			<=			16'h0101;
		end
		32'h0000C260: begin
				q			<=			16'h8067;
		end
		32'h0000C262: begin
				q			<=			16'h0000;
		end
		32'h0000C264: begin
				q			<=			16'h9863;
		end
		32'h0000C266: begin
				q			<=			16'h02A6;
		end
		32'h0000C268: begin
				q			<=			16'hEFB3;
		end
		32'h0000C26A: begin
				q			<=			16'h0062;
		end
		32'h0000C26C: begin
				q			<=			16'hEFB3;
		end
		32'h0000C26E: begin
				q			<=			16'h01CF;
		end
		32'h0000C270: begin
				q			<=			16'hEFB3;
		end
		32'h0000C272: begin
				q			<=			16'h01DF;
		end
		32'h0000C274: begin
				q			<=			16'h0513;
		end
		32'h0000C276: begin
				q			<=			16'h0020;
		end
		32'h0000C278: begin
				q			<=			16'h92E3;
		end
		32'h0000C27A: begin
				q			<=			16'hFE0F;
		end
		32'h0000C27C: begin
				q			<=			16'h1263;
		end
		32'h0000C27E: begin
				q			<=			16'h0407;
		end
		32'h0000C280: begin
				q			<=			16'h6533;
		end
		32'h0000C282: begin
				q			<=			16'h00CF;
		end
		32'h0000C284: begin
				q			<=			16'h6533;
		end
		32'h0000C286: begin
				q			<=			16'h0105;
		end
		32'h0000C288: begin
				q			<=			16'h6533;
		end
		32'h0000C28A: begin
				q			<=			16'h00B5;
		end
		32'h0000C28C: begin
				q			<=			16'h3513;
		end
		32'h0000C28E: begin
				q			<=			16'h0015;
		end
		32'h0000C290: begin
				q			<=			16'h006F;
		end
		32'h0000C292: begin
				q			<=			16'h02C0;
		end
		32'h0000C294: begin
				q			<=			16'h1463;
		end
		32'h0000C296: begin
				q			<=			16'h0A07;
		end
		32'h0000C298: begin
				q			<=			16'h6533;
		end
		32'h0000C29A: begin
				q			<=			16'h00CF;
		end
		32'h0000C29C: begin
				q			<=			16'h6533;
		end
		32'h0000C29E: begin
				q			<=			16'h0105;
		end
		32'h0000C2A0: begin
				q			<=			16'h6533;
		end
		32'h0000C2A2: begin
				q			<=			16'h00B5;
		end
		32'h0000C2A4: begin
				q			<=			16'h3513;
		end
		32'h0000C2A6: begin
				q			<=			16'h0015;
		end
		32'h0000C2A8: begin
				q			<=			16'h9A63;
		end
		32'h0000C2AA: begin
				q			<=			16'h0006;
		end
		32'h0000C2AC: begin
				q			<=			16'hEFB3;
		end
		32'h0000C2AE: begin
				q			<=			16'h0062;
		end
		32'h0000C2B0: begin
				q			<=			16'hEFB3;
		end
		32'h0000C2B2: begin
				q			<=			16'h01CF;
		end
		32'h0000C2B4: begin
				q			<=			16'hEFB3;
		end
		32'h0000C2B6: begin
				q			<=			16'h01DF;
		end
		32'h0000C2B8: begin
				q			<=			16'h8C63;
		end
		32'h0000C2BA: begin
				q			<=			16'h060F;
		end
		32'h0000C2BC: begin
				q			<=			16'h1A63;
		end
		32'h0000C2BE: begin
				q			<=			16'h0005;
		end
		32'h0000C2C0: begin
				q			<=			16'h8E63;
		end
		32'h0000C2C2: begin
				q			<=			16'h0117;
		end
		32'h0000C2C4: begin
				q			<=			16'h0513;
		end
		32'h0000C2C6: begin
				q			<=			16'h0010;
		end
		32'h0000C2C8: begin
				q			<=			16'h8AE3;
		end
		32'h0000C2CA: begin
				q			<=			16'hF807;
		end
		32'h0000C2CC: begin
				q			<=			16'h006F;
		end
		32'h0000C2CE: begin
				q			<=			16'h0080;
		end
		32'h0000C2D0: begin
				q			<=			16'h96E3;
		end
		32'h0000C2D2: begin
				q			<=			16'hF808;
		end
		32'h0000C2D4: begin
				q			<=			16'h0513;
		end
		32'h0000C2D6: begin
				q			<=			16'hFFF0;
		end
		32'h0000C2D8: begin
				q			<=			16'hF06F;
		end
		32'h0000C2DA: begin
				q			<=			16'hF85F;
		end
		32'h0000C2DC: begin
				q			<=			16'hC4E3;
		end
		32'h0000C2DE: begin
				q			<=			16'hFEE6;
		end
		32'h0000C2E0: begin
				q			<=			16'h5A63;
		end
		32'h0000C2E2: begin
				q			<=			16'h00D7;
		end
		32'h0000C2E4: begin
				q			<=			16'h0513;
		end
		32'h0000C2E6: begin
				q			<=			16'hFFF0;
		end
		32'h0000C2E8: begin
				q			<=			16'h8AE3;
		end
		32'h0000C2EA: begin
				q			<=			16'hF607;
		end
		32'h0000C2EC: begin
				q			<=			16'h0513;
		end
		32'h0000C2EE: begin
				q			<=			16'h0010;
		end
		32'h0000C2F0: begin
				q			<=			16'hF06F;
		end
		32'h0000C2F2: begin
				q			<=			16'hF6DF;
		end
		32'h0000C2F4: begin
				q			<=			16'hE8E3;
		end
		32'h0000C2F6: begin
				q			<=			16'hFCBE;
		end
		32'h0000C2F8: begin
				q			<=			16'h9663;
		end
		32'h0000C2FA: begin
				q			<=			16'h03D5;
		end
		32'h0000C2FC: begin
				q			<=			16'h64E3;
		end
		32'h0000C2FE: begin
				q			<=			16'hFD0E;
		end
		32'h0000C300: begin
				q			<=			16'h1463;
		end
		32'h0000C302: begin
				q			<=			16'h05C8;
		end
		32'h0000C304: begin
				q			<=			16'h60E3;
		end
		32'h0000C306: begin
				q			<=			16'hFCC3;
		end
		32'h0000C308: begin
				q			<=			16'h1463;
		end
		32'h0000C30A: begin
				q			<=			16'h0066;
		end
		32'h0000C30C: begin
				q			<=			16'hECE3;
		end
		32'h0000C30E: begin
				q			<=			16'hFBE2;
		end
		32'h0000C310: begin
				q			<=			16'h6AE3;
		end
		32'h0000C312: begin
				q			<=			16'hFC66;
		end
		32'h0000C314: begin
				q			<=			16'h0513;
		end
		32'h0000C316: begin
				q			<=			16'h0000;
		end
		32'h0000C318: begin
				q			<=			16'h12E3;
		end
		32'h0000C31A: begin
				q			<=			16'hF466;
		end
		32'h0000C31C: begin
				q			<=			16'h64E3;
		end
		32'h0000C31E: begin
				q			<=			16'hFC5F;
		end
		32'h0000C320: begin
				q			<=			16'hF06F;
		end
		32'h0000C322: begin
				q			<=			16'hF3DF;
		end
		32'h0000C324: begin
				q			<=			16'hE0E3;
		end
		32'h0000C326: begin
				q			<=			16'hFDD5;
		end
		32'h0000C328: begin
				q			<=			16'h0513;
		end
		32'h0000C32A: begin
				q			<=			16'h0000;
		end
		32'h0000C32C: begin
				q			<=			16'hF06F;
		end
		32'h0000C32E: begin
				q			<=			16'hF31F;
		end
		32'h0000C330: begin
				q			<=			16'h1CE3;
		end
		32'h0000C332: begin
				q			<=			16'hFE05;
		end
		32'h0000C334: begin
				q			<=			16'hF06F;
		end
		32'h0000C336: begin
				q			<=			16'hF91F;
		end
		32'h0000C338: begin
				q			<=			16'h88E3;
		end
		32'h0000C33A: begin
				q			<=			16'hF2E6;
		end
		32'h0000C33C: begin
				q			<=			16'h0513;
		end
		32'h0000C33E: begin
				q			<=			16'h0000;
		end
		32'h0000C340: begin
				q			<=			16'h86E3;
		end
		32'h0000C342: begin
				q			<=			16'hF606;
		end
		32'h0000C344: begin
				q			<=			16'hF06F;
		end
		32'h0000C346: begin
				q			<=			16'hF7DF;
		end
		32'h0000C348: begin
				q			<=			16'h6EE3;
		end
		32'h0000C34A: begin
				q			<=			16'hF9C8;
		end
		32'h0000C34C: begin
				q			<=			16'hF06F;
		end
		32'h0000C34E: begin
				q			<=			16'hFDDF;
		end
		32'h0000C350: begin
				q			<=			16'h0000;
		end
		32'h0000C352: begin
				q			<=			16'h0000;
		end
		32'h0000C354: begin
				q			<=			16'h0113;
		end
		32'h0000C356: begin
				q			<=			16'hF401;
		end
		32'h0000C358: begin
				q			<=			16'h2623;
		end
		32'h0000C35A: begin
				q			<=			16'h0B31;
		end
		32'h0000C35C: begin
				q			<=			16'hA983;
		end
		32'h0000C35E: begin
				q			<=			16'h00C5;
		end
		32'h0000C360: begin
				q			<=			16'hA683;
		end
		32'h0000C362: begin
				q			<=			16'h0005;
		end
		32'h0000C364: begin
				q			<=			16'hA783;
		end
		32'h0000C366: begin
				q			<=			16'h0045;
		end
		32'h0000C368: begin
				q			<=			16'h2623;
		end
		32'h0000C36A: begin
				q			<=			16'h00A1;
		end
		32'h0000C36C: begin
				q			<=			16'hA503;
		end
		32'h0000C36E: begin
				q			<=			16'h0085;
		end
		32'h0000C370: begin
				q			<=			16'h9713;
		end
		32'h0000C372: begin
				q			<=			16'h0109;
		end
		32'h0000C374: begin
				q			<=			16'h2823;
		end
		32'h0000C376: begin
				q			<=			16'h0B21;
		end
		32'h0000C378: begin
				q			<=			16'h2423;
		end
		32'h0000C37A: begin
				q			<=			16'h0B41;
		end
		32'h0000C37C: begin
				q			<=			16'h2223;
		end
		32'h0000C37E: begin
				q			<=			16'h0B51;
		end
		32'h0000C380: begin
				q			<=			16'h2023;
		end
		32'h0000C382: begin
				q			<=			16'h0B61;
		end
		32'h0000C384: begin
				q			<=			16'h2A03;
		end
		32'h0000C386: begin
				q			<=			16'h0006;
		end
		32'h0000C388: begin
				q			<=			16'h2B03;
		end
		32'h0000C38A: begin
				q			<=			16'h0046;
		end
		32'h0000C38C: begin
				q			<=			16'h2A83;
		end
		32'h0000C38E: begin
				q			<=			16'h0086;
		end
		32'h0000C390: begin
				q			<=			16'h2903;
		end
		32'h0000C392: begin
				q			<=			16'h00C6;
		end
		32'h0000C394: begin
				q			<=			16'h8637;
		end
		32'h0000C396: begin
				q			<=			16'h0000;
		end
		32'h0000C398: begin
				q			<=			16'h2A23;
		end
		32'h0000C39A: begin
				q			<=			16'h0A91;
		end
		32'h0000C39C: begin
				q			<=			16'h5713;
		end
		32'h0000C39E: begin
				q			<=			16'h0107;
		end
		32'h0000C3A0: begin
				q			<=			16'hD493;
		end
		32'h0000C3A2: begin
				q			<=			16'h0109;
		end
		32'h0000C3A4: begin
				q			<=			16'h0613;
		end
		32'h0000C3A6: begin
				q			<=			16'hFFF6;
		end
		32'h0000C3A8: begin
				q			<=			16'h2623;
		end
		32'h0000C3AA: begin
				q			<=			16'h0731;
		end
		32'h0000C3AC: begin
				q			<=			16'h2E23;
		end
		32'h0000C3AE: begin
				q			<=			16'h0A11;
		end
		32'h0000C3B0: begin
				q			<=			16'h2C23;
		end
		32'h0000C3B2: begin
				q			<=			16'h0A81;
		end
		32'h0000C3B4: begin
				q			<=			16'h2E23;
		end
		32'h0000C3B6: begin
				q			<=			16'h0971;
		end
		32'h0000C3B8: begin
				q			<=			16'h2C23;
		end
		32'h0000C3BA: begin
				q			<=			16'h0981;
		end
		32'h0000C3BC: begin
				q			<=			16'h2A23;
		end
		32'h0000C3BE: begin
				q			<=			16'h0991;
		end
		32'h0000C3C0: begin
				q			<=			16'h2823;
		end
		32'h0000C3C2: begin
				q			<=			16'h09A1;
		end
		32'h0000C3C4: begin
				q			<=			16'h2623;
		end
		32'h0000C3C6: begin
				q			<=			16'h09B1;
		end
		32'h0000C3C8: begin
				q			<=			16'h2023;
		end
		32'h0000C3CA: begin
				q			<=			16'h06D1;
		end
		32'h0000C3CC: begin
				q			<=			16'h2223;
		end
		32'h0000C3CE: begin
				q			<=			16'h06F1;
		end
		32'h0000C3D0: begin
				q			<=			16'h2423;
		end
		32'h0000C3D2: begin
				q			<=			16'h06A1;
		end
		32'h0000C3D4: begin
				q			<=			16'h2823;
		end
		32'h0000C3D6: begin
				q			<=			16'h02D1;
		end
		32'h0000C3D8: begin
				q			<=			16'h2A23;
		end
		32'h0000C3DA: begin
				q			<=			16'h02F1;
		end
		32'h0000C3DC: begin
				q			<=			16'h2C23;
		end
		32'h0000C3DE: begin
				q			<=			16'h02A1;
		end
		32'h0000C3E0: begin
				q			<=			16'h2E23;
		end
		32'h0000C3E2: begin
				q			<=			16'h02E1;
		end
		32'h0000C3E4: begin
				q			<=			16'h74B3;
		end
		32'h0000C3E6: begin
				q			<=			16'h0096;
		end
		32'h0000C3E8: begin
				q			<=			16'hD993;
		end
		32'h0000C3EA: begin
				q			<=			16'h01F9;
		end
		32'h0000C3EC: begin
				q			<=			16'h8A63;
		end
		32'h0000C3EE: begin
				q			<=			16'h1204;
		end
		32'h0000C3F0: begin
				q			<=			16'h8A63;
		end
		32'h0000C3F2: begin
				q			<=			16'h24C4;
		end
		32'h0000C3F4: begin
				q			<=			16'h07B7;
		end
		32'h0000C3F6: begin
				q			<=			16'h0001;
		end
		32'h0000C3F8: begin
				q			<=			16'h67B3;
		end
		32'h0000C3FA: begin
				q			<=			16'h00F7;
		end
		32'h0000C3FC: begin
				q			<=			16'h2E23;
		end
		32'h0000C3FE: begin
				q			<=			16'h02F1;
		end
		32'h0000C400: begin
				q			<=			16'h0613;
		end
		32'h0000C402: begin
				q			<=			16'h0301;
		end
		32'h0000C404: begin
				q			<=			16'h0793;
		end
		32'h0000C406: begin
				q			<=			16'h03C1;
		end
		32'h0000C408: begin
				q			<=			16'hA703;
		end
		32'h0000C40A: begin
				q			<=			16'h0007;
		end
		32'h0000C40C: begin
				q			<=			16'hA683;
		end
		32'h0000C40E: begin
				q			<=			16'hFFC7;
		end
		32'h0000C410: begin
				q			<=			16'h8793;
		end
		32'h0000C412: begin
				q			<=			16'hFFC7;
		end
		32'h0000C414: begin
				q			<=			16'h1713;
		end
		32'h0000C416: begin
				q			<=			16'h0037;
		end
		32'h0000C418: begin
				q			<=			16'hD693;
		end
		32'h0000C41A: begin
				q			<=			16'h01D6;
		end
		32'h0000C41C: begin
				q			<=			16'h6733;
		end
		32'h0000C41E: begin
				q			<=			16'h00D7;
		end
		32'h0000C420: begin
				q			<=			16'hA223;
		end
		32'h0000C422: begin
				q			<=			16'h00E7;
		end
		32'h0000C424: begin
				q			<=			16'h12E3;
		end
		32'h0000C426: begin
				q			<=			16'hFEF6;
		end
		32'h0000C428: begin
				q			<=			16'h2783;
		end
		32'h0000C42A: begin
				q			<=			16'h0301;
		end
		32'h0000C42C: begin
				q			<=			16'hC537;
		end
		32'h0000C42E: begin
				q			<=			16'hFFFF;
		end
		32'h0000C430: begin
				q			<=			16'h0513;
		end
		32'h0000C432: begin
				q			<=			16'h0015;
		end
		32'h0000C434: begin
				q			<=			16'h9793;
		end
		32'h0000C436: begin
				q			<=			16'h0037;
		end
		32'h0000C438: begin
				q			<=			16'h2823;
		end
		32'h0000C43A: begin
				q			<=			16'h02F1;
		end
		32'h0000C43C: begin
				q			<=			16'h84B3;
		end
		32'h0000C43E: begin
				q			<=			16'h00A4;
		end
		32'h0000C440: begin
				q			<=			16'h0B93;
		end
		32'h0000C442: begin
				q			<=			16'h0000;
		end
		32'h0000C444: begin
				q			<=			16'h1793;
		end
		32'h0000C446: begin
				q			<=			16'h0109;
		end
		32'h0000C448: begin
				q			<=			16'h8737;
		end
		32'h0000C44A: begin
				q			<=			16'h0000;
		end
		32'h0000C44C: begin
				q			<=			16'h5513;
		end
		32'h0000C44E: begin
				q			<=			16'h0109;
		end
		32'h0000C450: begin
				q			<=			16'hD793;
		end
		32'h0000C452: begin
				q			<=			16'h0107;
		end
		32'h0000C454: begin
				q			<=			16'h0713;
		end
		32'h0000C456: begin
				q			<=			16'hFFF7;
		end
		32'h0000C458: begin
				q			<=			16'h2623;
		end
		32'h0000C45A: begin
				q			<=			16'h0721;
		end
		32'h0000C45C: begin
				q			<=			16'h2023;
		end
		32'h0000C45E: begin
				q			<=			16'h0741;
		end
		32'h0000C460: begin
				q			<=			16'h2223;
		end
		32'h0000C462: begin
				q			<=			16'h0761;
		end
		32'h0000C464: begin
				q			<=			16'h2423;
		end
		32'h0000C466: begin
				q			<=			16'h0751;
		end
		32'h0000C468: begin
				q			<=			16'h2023;
		end
		32'h0000C46A: begin
				q			<=			16'h0541;
		end
		32'h0000C46C: begin
				q			<=			16'h2223;
		end
		32'h0000C46E: begin
				q			<=			16'h0561;
		end
		32'h0000C470: begin
				q			<=			16'h2423;
		end
		32'h0000C472: begin
				q			<=			16'h0551;
		end
		32'h0000C474: begin
				q			<=			16'h2623;
		end
		32'h0000C476: begin
				q			<=			16'h04F1;
		end
		32'h0000C478: begin
				q			<=			16'h7533;
		end
		32'h0000C47A: begin
				q			<=			16'h00A7;
		end
		32'h0000C47C: begin
				q			<=			16'h5913;
		end
		32'h0000C47E: begin
				q			<=			16'h01F9;
		end
		32'h0000C480: begin
				q			<=			16'h0663;
		end
		32'h0000C482: begin
				q			<=			16'h1E05;
		end
		32'h0000C484: begin
				q			<=			16'h0863;
		end
		32'h0000C486: begin
				q			<=			16'h30E5;
		end
		32'h0000C488: begin
				q			<=			16'h0AB7;
		end
		32'h0000C48A: begin
				q			<=			16'h0001;
		end
		32'h0000C48C: begin
				q			<=			16'hEAB3;
		end
		32'h0000C48E: begin
				q			<=			16'h0157;
		end
		32'h0000C490: begin
				q			<=			16'h2623;
		end
		32'h0000C492: begin
				q			<=			16'h0551;
		end
		32'h0000C494: begin
				q			<=			16'h0613;
		end
		32'h0000C496: begin
				q			<=			16'h0401;
		end
		32'h0000C498: begin
				q			<=			16'h0793;
		end
		32'h0000C49A: begin
				q			<=			16'h04C1;
		end
		32'h0000C49C: begin
				q			<=			16'hA703;
		end
		32'h0000C49E: begin
				q			<=			16'h0007;
		end
		32'h0000C4A0: begin
				q			<=			16'hA683;
		end
		32'h0000C4A2: begin
				q			<=			16'hFFC7;
		end
		32'h0000C4A4: begin
				q			<=			16'h8793;
		end
		32'h0000C4A6: begin
				q			<=			16'hFFC7;
		end
		32'h0000C4A8: begin
				q			<=			16'h1713;
		end
		32'h0000C4AA: begin
				q			<=			16'h0037;
		end
		32'h0000C4AC: begin
				q			<=			16'hD693;
		end
		32'h0000C4AE: begin
				q			<=			16'h01D6;
		end
		32'h0000C4B0: begin
				q			<=			16'h6733;
		end
		32'h0000C4B2: begin
				q			<=			16'h00D7;
		end
		32'h0000C4B4: begin
				q			<=			16'hA223;
		end
		32'h0000C4B6: begin
				q			<=			16'h00E7;
		end
		32'h0000C4B8: begin
				q			<=			16'h12E3;
		end
		32'h0000C4BA: begin
				q			<=			16'hFEF6;
		end
		32'h0000C4BC: begin
				q			<=			16'h2783;
		end
		32'h0000C4BE: begin
				q			<=			16'h0401;
		end
		32'h0000C4C0: begin
				q			<=			16'h9793;
		end
		32'h0000C4C2: begin
				q			<=			16'h0037;
		end
		32'h0000C4C4: begin
				q			<=			16'h2023;
		end
		32'h0000C4C6: begin
				q			<=			16'h04F1;
		end
		32'h0000C4C8: begin
				q			<=			16'hC7B7;
		end
		32'h0000C4CA: begin
				q			<=			16'hFFFF;
		end
		32'h0000C4CC: begin
				q			<=			16'h8793;
		end
		32'h0000C4CE: begin
				q			<=			16'h0017;
		end
		32'h0000C4D0: begin
				q			<=			16'h0533;
		end
		32'h0000C4D2: begin
				q			<=			16'h00F5;
		end
		32'h0000C4D4: begin
				q			<=			16'h0713;
		end
		32'h0000C4D6: begin
				q			<=			16'h0000;
		end
		32'h0000C4D8: begin
				q			<=			16'hC7B3;
		end
		32'h0000C4DA: begin
				q			<=			16'h0129;
		end
		32'h0000C4DC: begin
				q			<=			16'h2823;
		end
		32'h0000C4DE: begin
				q			<=			16'h00F1;
		end
		32'h0000C4E0: begin
				q			<=			16'h07B3;
		end
		32'h0000C4E2: begin
				q			<=			16'h0095;
		end
		32'h0000C4E4: begin
				q			<=			16'h2023;
		end
		32'h0000C4E6: begin
				q			<=			16'h02F1;
		end
		32'h0000C4E8: begin
				q			<=			16'h8793;
		end
		32'h0000C4EA: begin
				q			<=			16'h0017;
		end
		32'h0000C4EC: begin
				q			<=			16'h2E23;
		end
		32'h0000C4EE: begin
				q			<=			16'h00F1;
		end
		32'h0000C4F0: begin
				q			<=			16'h9793;
		end
		32'h0000C4F2: begin
				q			<=			16'h002B;
		end
		32'h0000C4F4: begin
				q			<=			16'hE7B3;
		end
		32'h0000C4F6: begin
				q			<=			16'h00E7;
		end
		32'h0000C4F8: begin
				q			<=			16'h8793;
		end
		32'h0000C4FA: begin
				q			<=			16'hFFF7;
		end
		32'h0000C4FC: begin
				q			<=			16'h0693;
		end
		32'h0000C4FE: begin
				q			<=			16'h00E0;
		end
		32'h0000C500: begin
				q			<=			16'hEE63;
		end
		32'h0000C502: begin
				q			<=			16'h2AF6;
		end
		32'h0000C504: begin
				q			<=			16'h3697;
		end
		32'h0000C506: begin
				q			<=			16'h0000;
		end
		32'h0000C508: begin
				q			<=			16'h8693;
		end
		32'h0000C50A: begin
				q			<=			16'h42C6;
		end
		32'h0000C50C: begin
				q			<=			16'h9793;
		end
		32'h0000C50E: begin
				q			<=			16'h0027;
		end
		32'h0000C510: begin
				q			<=			16'h87B3;
		end
		32'h0000C512: begin
				q			<=			16'h00D7;
		end
		32'h0000C514: begin
				q			<=			16'hA783;
		end
		32'h0000C516: begin
				q			<=			16'h0007;
		end
		32'h0000C518: begin
				q			<=			16'h87B3;
		end
		32'h0000C51A: begin
				q			<=			16'h00D7;
		end
		32'h0000C51C: begin
				q			<=			16'h8067;
		end
		32'h0000C51E: begin
				q			<=			16'h0007;
		end
		32'h0000C520: begin
				q			<=			16'hE633;
		end
		32'h0000C522: begin
				q			<=			16'h00D7;
		end
		32'h0000C524: begin
				q			<=			16'h6633;
		end
		32'h0000C526: begin
				q			<=			16'h00A6;
		end
		32'h0000C528: begin
				q			<=			16'h6633;
		end
		32'h0000C52A: begin
				q			<=			16'h00E6;
		end
		32'h0000C52C: begin
				q			<=			16'h0A63;
		end
		32'h0000C52E: begin
				q			<=			16'h1206;
		end
		32'h0000C530: begin
				q			<=			16'h0C63;
		end
		32'h0000C532: begin
				q			<=			16'h0407;
		end
		32'h0000C534: begin
				q			<=			16'h0513;
		end
		32'h0000C536: begin
				q			<=			16'h0007;
		end
		32'h0000C538: begin
				q			<=			16'h20EF;
		end
		32'h0000C53A: begin
				q			<=			16'h3950;
		end
		32'h0000C53C: begin
				q			<=			16'h0713;
		end
		32'h0000C53E: begin
				q			<=			16'hFF45;
		end
		32'h0000C540: begin
				q			<=			16'h5793;
		end
		32'h0000C542: begin
				q			<=			16'h4057;
		end
		32'h0000C544: begin
				q			<=			16'h7713;
		end
		32'h0000C546: begin
				q			<=			16'h01F7;
		end
		32'h0000C548: begin
				q			<=			16'h0A63;
		end
		32'h0000C54A: begin
				q			<=			16'h0607;
		end
		32'h0000C54C: begin
				q			<=			16'h0693;
		end
		32'h0000C54E: begin
				q			<=			16'hFFC0;
		end
		32'h0000C550: begin
				q			<=			16'h86B3;
		end
		32'h0000C552: begin
				q			<=			16'h02D7;
		end
		32'h0000C554: begin
				q			<=			16'h0813;
		end
		32'h0000C556: begin
				q			<=			16'h0200;
		end
		32'h0000C558: begin
				q			<=			16'h9593;
		end
		32'h0000C55A: begin
				q			<=			16'h0027;
		end
		32'h0000C55C: begin
				q			<=			16'h0E13;
		end
		32'h0000C55E: begin
				q			<=			16'hFF00;
		end
		32'h0000C560: begin
				q			<=			16'h0833;
		end
		32'h0000C562: begin
				q			<=			16'h40E8;
		end
		32'h0000C564: begin
				q			<=			16'h8693;
		end
		32'h0000C566: begin
				q			<=			16'hFFC6;
		end
		32'h0000C568: begin
				q			<=			16'h9C63;
		end
		32'h0000C56A: begin
				q			<=			16'h09C6;
		end
		32'h0000C56C: begin
				q			<=			16'h0693;
		end
		32'h0000C56E: begin
				q			<=			16'h0801;
		end
		32'h0000C570: begin
				q			<=			16'h85B3;
		end
		32'h0000C572: begin
				q			<=			16'h00B6;
		end
		32'h0000C574: begin
				q			<=			16'h2683;
		end
		32'h0000C576: begin
				q			<=			16'h0301;
		end
		32'h0000C578: begin
				q			<=			16'h8793;
		end
		32'h0000C57A: begin
				q			<=			16'hFFF7;
		end
		32'h0000C57C: begin
				q			<=			16'h9733;
		end
		32'h0000C57E: begin
				q			<=			16'h00E6;
		end
		32'h0000C580: begin
				q			<=			16'hA823;
		end
		32'h0000C582: begin
				q			<=			16'hFAE5;
		end
		32'h0000C584: begin
				q			<=			16'h006F;
		end
		32'h0000C586: begin
				q			<=			16'h0640;
		end
		32'h0000C588: begin
				q			<=			16'h0863;
		end
		32'h0000C58A: begin
				q			<=			16'h0005;
		end
		32'h0000C58C: begin
				q			<=			16'h20EF;
		end
		32'h0000C58E: begin
				q			<=			16'h3410;
		end
		32'h0000C590: begin
				q			<=			16'h0513;
		end
		32'h0000C592: begin
				q			<=			16'h0205;
		end
		32'h0000C594: begin
				q			<=			16'hF06F;
		end
		32'h0000C596: begin
				q			<=			16'hFA9F;
		end
		32'h0000C598: begin
				q			<=			16'h8A63;
		end
		32'h0000C59A: begin
				q			<=			16'h0007;
		end
		32'h0000C59C: begin
				q			<=			16'h8513;
		end
		32'h0000C59E: begin
				q			<=			16'h0007;
		end
		32'h0000C5A0: begin
				q			<=			16'h20EF;
		end
		32'h0000C5A2: begin
				q			<=			16'h32D0;
		end
		32'h0000C5A4: begin
				q			<=			16'h0513;
		end
		32'h0000C5A6: begin
				q			<=			16'h0405;
		end
		32'h0000C5A8: begin
				q			<=			16'hF06F;
		end
		32'h0000C5AA: begin
				q			<=			16'hF95F;
		end
		32'h0000C5AC: begin
				q			<=			16'h8513;
		end
		32'h0000C5AE: begin
				q			<=			16'h0006;
		end
		32'h0000C5B0: begin
				q			<=			16'h20EF;
		end
		32'h0000C5B2: begin
				q			<=			16'h31D0;
		end
		32'h0000C5B4: begin
				q			<=			16'h0513;
		end
		32'h0000C5B6: begin
				q			<=			16'h0605;
		end
		32'h0000C5B8: begin
				q			<=			16'hF06F;
		end
		32'h0000C5BA: begin
				q			<=			16'hF85F;
		end
		32'h0000C5BC: begin
				q			<=			16'h0613;
		end
		32'h0000C5BE: begin
				q			<=			16'hFFC0;
		end
		32'h0000C5C0: begin
				q			<=			16'h8633;
		end
		32'h0000C5C2: begin
				q			<=			16'h02C7;
		end
		32'h0000C5C4: begin
				q			<=			16'h0713;
		end
		32'h0000C5C6: begin
				q			<=			16'h0301;
		end
		32'h0000C5C8: begin
				q			<=			16'h0693;
		end
		32'h0000C5CA: begin
				q			<=			16'h0030;
		end
		32'h0000C5CC: begin
				q			<=			16'h05B3;
		end
		32'h0000C5CE: begin
				q			<=			16'h00C7;
		end
		32'h0000C5D0: begin
				q			<=			16'hA583;
		end
		32'h0000C5D2: begin
				q			<=			16'h00C5;
		end
		32'h0000C5D4: begin
				q			<=			16'h8693;
		end
		32'h0000C5D6: begin
				q			<=			16'hFFF6;
		end
		32'h0000C5D8: begin
				q			<=			16'h0713;
		end
		32'h0000C5DA: begin
				q			<=			16'hFFC7;
		end
		32'h0000C5DC: begin
				q			<=			16'h2823;
		end
		32'h0000C5DE: begin
				q			<=			16'h00B7;
		end
		32'h0000C5E0: begin
				q			<=			16'hD6E3;
		end
		32'h0000C5E2: begin
				q			<=			16'hFEF6;
		end
		32'h0000C5E4: begin
				q			<=			16'h8793;
		end
		32'h0000C5E6: begin
				q			<=			16'hFFF7;
		end
		32'h0000C5E8: begin
				q			<=			16'h0693;
		end
		32'h0000C5EA: begin
				q			<=			16'hFFF0;
		end
		32'h0000C5EC: begin
				q			<=			16'h9063;
		end
		32'h0000C5EE: begin
				q			<=			16'h04D7;
		end
		32'h0000C5F0: begin
				q			<=			16'hC4B7;
		end
		32'h0000C5F2: begin
				q			<=			16'hFFFF;
		end
		32'h0000C5F4: begin
				q			<=			16'h8493;
		end
		32'h0000C5F6: begin
				q			<=			16'h0114;
		end
		32'h0000C5F8: begin
				q			<=			16'h84B3;
		end
		32'h0000C5FA: begin
				q			<=			16'h40A4;
		end
		32'h0000C5FC: begin
				q			<=			16'hF06F;
		end
		32'h0000C5FE: begin
				q			<=			16'hE45F;
		end
		32'h0000C600: begin
				q			<=			16'h0613;
		end
		32'h0000C602: begin
				q			<=			16'h0301;
		end
		32'h0000C604: begin
				q			<=			16'h0333;
		end
		32'h0000C606: begin
				q			<=			16'h00D6;
		end
		32'h0000C608: begin
				q			<=			16'h88B3;
		end
		32'h0000C60A: begin
				q			<=			16'h00D5;
		end
		32'h0000C60C: begin
				q			<=			16'h08B3;
		end
		32'h0000C60E: begin
				q			<=			16'h0116;
		end
		32'h0000C610: begin
				q			<=			16'h2603;
		end
		32'h0000C612: begin
				q			<=			16'h00C3;
		end
		32'h0000C614: begin
				q			<=			16'h2303;
		end
		32'h0000C616: begin
				q			<=			16'h0103;
		end
		32'h0000C618: begin
				q			<=			16'h5633;
		end
		32'h0000C61A: begin
				q			<=			16'h0106;
		end
		32'h0000C61C: begin
				q			<=			16'h1333;
		end
		32'h0000C61E: begin
				q			<=			16'h00E3;
		end
		32'h0000C620: begin
				q			<=			16'h6633;
		end
		32'h0000C622: begin
				q			<=			16'h0066;
		end
		32'h0000C624: begin
				q			<=			16'hA823;
		end
		32'h0000C626: begin
				q			<=			16'h00C8;
		end
		32'h0000C628: begin
				q			<=			16'hF06F;
		end
		32'h0000C62A: begin
				q			<=			16'hF3DF;
		end
		32'h0000C62C: begin
				q			<=			16'h9713;
		end
		32'h0000C62E: begin
				q			<=			16'h0027;
		end
		32'h0000C630: begin
				q			<=			16'h0613;
		end
		32'h0000C632: begin
				q			<=			16'h0301;
		end
		32'h0000C634: begin
				q			<=			16'h0733;
		end
		32'h0000C636: begin
				q			<=			16'h00E6;
		end
		32'h0000C638: begin
				q			<=			16'h2023;
		end
		32'h0000C63A: begin
				q			<=			16'h0007;
		end
		32'h0000C63C: begin
				q			<=			16'h8793;
		end
		32'h0000C63E: begin
				q			<=			16'hFFF7;
		end
		32'h0000C640: begin
				q			<=			16'hF06F;
		end
		32'h0000C642: begin
				q			<=			16'hFADF;
		end
		32'h0000C644: begin
				q			<=			16'hE7B3;
		end
		32'h0000C646: begin
				q			<=			16'h00D7;
		end
		32'h0000C648: begin
				q			<=			16'hE7B3;
		end
		32'h0000C64A: begin
				q			<=			16'h00A7;
		end
		32'h0000C64C: begin
				q			<=			16'hE7B3;
		end
		32'h0000C64E: begin
				q			<=			16'h00E7;
		end
		32'h0000C650: begin
				q			<=			16'h0B93;
		end
		32'h0000C652: begin
				q			<=			16'h0020;
		end
		32'h0000C654: begin
				q			<=			16'h88E3;
		end
		32'h0000C656: begin
				q			<=			16'hDE07;
		end
		32'h0000C658: begin
				q			<=			16'h0B93;
		end
		32'h0000C65A: begin
				q			<=			16'h0030;
		end
		32'h0000C65C: begin
				q			<=			16'hF06F;
		end
		32'h0000C65E: begin
				q			<=			16'hDE9F;
		end
		32'h0000C660: begin
				q			<=			16'h0493;
		end
		32'h0000C662: begin
				q			<=			16'h0000;
		end
		32'h0000C664: begin
				q			<=			16'h0B93;
		end
		32'h0000C666: begin
				q			<=			16'h0010;
		end
		32'h0000C668: begin
				q			<=			16'hF06F;
		end
		32'h0000C66A: begin
				q			<=			16'hDDDF;
		end
		32'h0000C66C: begin
				q			<=			16'h6733;
		end
		32'h0000C66E: begin
				q			<=			16'h016A;
		end
		32'h0000C670: begin
				q			<=			16'h6733;
		end
		32'h0000C672: begin
				q			<=			16'h0157;
		end
		32'h0000C674: begin
				q			<=			16'h6733;
		end
		32'h0000C676: begin
				q			<=			16'h00F7;
		end
		32'h0000C678: begin
				q			<=			16'h0C63;
		end
		32'h0000C67A: begin
				q			<=			16'h1207;
		end
		32'h0000C67C: begin
				q			<=			16'h8C63;
		end
		32'h0000C67E: begin
				q			<=			16'h0407;
		end
		32'h0000C680: begin
				q			<=			16'h8513;
		end
		32'h0000C682: begin
				q			<=			16'h0007;
		end
		32'h0000C684: begin
				q			<=			16'h20EF;
		end
		32'h0000C686: begin
				q			<=			16'h2490;
		end
		32'h0000C688: begin
				q			<=			16'h0713;
		end
		32'h0000C68A: begin
				q			<=			16'hFF45;
		end
		32'h0000C68C: begin
				q			<=			16'h5793;
		end
		32'h0000C68E: begin
				q			<=			16'h4057;
		end
		32'h0000C690: begin
				q			<=			16'h7713;
		end
		32'h0000C692: begin
				q			<=			16'h01F7;
		end
		32'h0000C694: begin
				q			<=			16'h0C63;
		end
		32'h0000C696: begin
				q			<=			16'h0607;
		end
		32'h0000C698: begin
				q			<=			16'h0693;
		end
		32'h0000C69A: begin
				q			<=			16'hFFC0;
		end
		32'h0000C69C: begin
				q			<=			16'h86B3;
		end
		32'h0000C69E: begin
				q			<=			16'h02D7;
		end
		32'h0000C6A0: begin
				q			<=			16'h0813;
		end
		32'h0000C6A2: begin
				q			<=			16'h0200;
		end
		32'h0000C6A4: begin
				q			<=			16'h9593;
		end
		32'h0000C6A6: begin
				q			<=			16'h0027;
		end
		32'h0000C6A8: begin
				q			<=			16'h0E13;
		end
		32'h0000C6AA: begin
				q			<=			16'hFF00;
		end
		32'h0000C6AC: begin
				q			<=			16'h0833;
		end
		32'h0000C6AE: begin
				q			<=			16'h40E8;
		end
		32'h0000C6B0: begin
				q			<=			16'h8693;
		end
		32'h0000C6B2: begin
				q			<=			16'hFFC6;
		end
		32'h0000C6B4: begin
				q			<=			16'h9E63;
		end
		32'h0000C6B6: begin
				q			<=			16'h09C6;
		end
		32'h0000C6B8: begin
				q			<=			16'h0693;
		end
		32'h0000C6BA: begin
				q			<=			16'h0801;
		end
		32'h0000C6BC: begin
				q			<=			16'h85B3;
		end
		32'h0000C6BE: begin
				q			<=			16'h00B6;
		end
		32'h0000C6C0: begin
				q			<=			16'h2683;
		end
		32'h0000C6C2: begin
				q			<=			16'h0401;
		end
		32'h0000C6C4: begin
				q			<=			16'h8793;
		end
		32'h0000C6C6: begin
				q			<=			16'hFFF7;
		end
		32'h0000C6C8: begin
				q			<=			16'h9733;
		end
		32'h0000C6CA: begin
				q			<=			16'h00E6;
		end
		32'h0000C6CC: begin
				q			<=			16'hA023;
		end
		32'h0000C6CE: begin
				q			<=			16'hFCE5;
		end
		32'h0000C6D0: begin
				q			<=			16'h006F;
		end
		32'h0000C6D2: begin
				q			<=			16'h0680;
		end
		32'h0000C6D4: begin
				q			<=			16'h8A63;
		end
		32'h0000C6D6: begin
				q			<=			16'h000A;
		end
		32'h0000C6D8: begin
				q			<=			16'h8513;
		end
		32'h0000C6DA: begin
				q			<=			16'h000A;
		end
		32'h0000C6DC: begin
				q			<=			16'h20EF;
		end
		32'h0000C6DE: begin
				q			<=			16'h1F10;
		end
		32'h0000C6E0: begin
				q			<=			16'h0513;
		end
		32'h0000C6E2: begin
				q			<=			16'h0205;
		end
		32'h0000C6E4: begin
				q			<=			16'hF06F;
		end
		32'h0000C6E6: begin
				q			<=			16'hFA5F;
		end
		32'h0000C6E8: begin
				q			<=			16'h0A63;
		end
		32'h0000C6EA: begin
				q			<=			16'h000B;
		end
		32'h0000C6EC: begin
				q			<=			16'h0513;
		end
		32'h0000C6EE: begin
				q			<=			16'h000B;
		end
		32'h0000C6F0: begin
				q			<=			16'h20EF;
		end
		32'h0000C6F2: begin
				q			<=			16'h1DD0;
		end
		32'h0000C6F4: begin
				q			<=			16'h0513;
		end
		32'h0000C6F6: begin
				q			<=			16'h0405;
		end
		32'h0000C6F8: begin
				q			<=			16'hF06F;
		end
		32'h0000C6FA: begin
				q			<=			16'hF91F;
		end
		32'h0000C6FC: begin
				q			<=			16'h0513;
		end
		32'h0000C6FE: begin
				q			<=			16'h000A;
		end
		32'h0000C700: begin
				q			<=			16'h20EF;
		end
		32'h0000C702: begin
				q			<=			16'h1CD0;
		end
		32'h0000C704: begin
				q			<=			16'h0513;
		end
		32'h0000C706: begin
				q			<=			16'h0605;
		end
		32'h0000C708: begin
				q			<=			16'hF06F;
		end
		32'h0000C70A: begin
				q			<=			16'hF81F;
		end
		32'h0000C70C: begin
				q			<=			16'h0613;
		end
		32'h0000C70E: begin
				q			<=			16'hFFC0;
		end
		32'h0000C710: begin
				q			<=			16'h8633;
		end
		32'h0000C712: begin
				q			<=			16'h02C7;
		end
		32'h0000C714: begin
				q			<=			16'h0713;
		end
		32'h0000C716: begin
				q			<=			16'h0401;
		end
		32'h0000C718: begin
				q			<=			16'h0693;
		end
		32'h0000C71A: begin
				q			<=			16'h0030;
		end
		32'h0000C71C: begin
				q			<=			16'h05B3;
		end
		32'h0000C71E: begin
				q			<=			16'h00C7;
		end
		32'h0000C720: begin
				q			<=			16'hA583;
		end
		32'h0000C722: begin
				q			<=			16'h00C5;
		end
		32'h0000C724: begin
				q			<=			16'h8693;
		end
		32'h0000C726: begin
				q			<=			16'hFFF6;
		end
		32'h0000C728: begin
				q			<=			16'h0713;
		end
		32'h0000C72A: begin
				q			<=			16'hFFC7;
		end
		32'h0000C72C: begin
				q			<=			16'h2823;
		end
		32'h0000C72E: begin
				q			<=			16'h00B7;
		end
		32'h0000C730: begin
				q			<=			16'hD6E3;
		end
		32'h0000C732: begin
				q			<=			16'hFEF6;
		end
		32'h0000C734: begin
				q			<=			16'h8793;
		end
		32'h0000C736: begin
				q			<=			16'hFFF7;
		end
		32'h0000C738: begin
				q			<=			16'h0693;
		end
		32'h0000C73A: begin
				q			<=			16'hFFF0;
		end
		32'h0000C73C: begin
				q			<=			16'h9063;
		end
		32'h0000C73E: begin
				q			<=			16'h04D7;
		end
		32'h0000C740: begin
				q			<=			16'hC7B7;
		end
		32'h0000C742: begin
				q			<=			16'hFFFF;
		end
		32'h0000C744: begin
				q			<=			16'h8793;
		end
		32'h0000C746: begin
				q			<=			16'h0117;
		end
		32'h0000C748: begin
				q			<=			16'h8533;
		end
		32'h0000C74A: begin
				q			<=			16'h40A7;
		end
		32'h0000C74C: begin
				q			<=			16'hF06F;
		end
		32'h0000C74E: begin
				q			<=			16'hD89F;
		end
		32'h0000C750: begin
				q			<=			16'h0613;
		end
		32'h0000C752: begin
				q			<=			16'h0401;
		end
		32'h0000C754: begin
				q			<=			16'h0333;
		end
		32'h0000C756: begin
				q			<=			16'h00D6;
		end
		32'h0000C758: begin
				q			<=			16'h88B3;
		end
		32'h0000C75A: begin
				q			<=			16'h00D5;
		end
		32'h0000C75C: begin
				q			<=			16'h08B3;
		end
		32'h0000C75E: begin
				q			<=			16'h0116;
		end
		32'h0000C760: begin
				q			<=			16'h2603;
		end
		32'h0000C762: begin
				q			<=			16'h00C3;
		end
		32'h0000C764: begin
				q			<=			16'h2303;
		end
		32'h0000C766: begin
				q			<=			16'h0103;
		end
		32'h0000C768: begin
				q			<=			16'h5633;
		end
		32'h0000C76A: begin
				q			<=			16'h0106;
		end
		32'h0000C76C: begin
				q			<=			16'h1333;
		end
		32'h0000C76E: begin
				q			<=			16'h00E3;
		end
		32'h0000C770: begin
				q			<=			16'h6633;
		end
		32'h0000C772: begin
				q			<=			16'h0066;
		end
		32'h0000C774: begin
				q			<=			16'hA823;
		end
		32'h0000C776: begin
				q			<=			16'h00C8;
		end
		32'h0000C778: begin
				q			<=			16'hF06F;
		end
		32'h0000C77A: begin
				q			<=			16'hF39F;
		end
		32'h0000C77C: begin
				q			<=			16'h9713;
		end
		32'h0000C77E: begin
				q			<=			16'h0027;
		end
		32'h0000C780: begin
				q			<=			16'h0613;
		end
		32'h0000C782: begin
				q			<=			16'h0401;
		end
		32'h0000C784: begin
				q			<=			16'h0733;
		end
		32'h0000C786: begin
				q			<=			16'h00E6;
		end
		32'h0000C788: begin
				q			<=			16'h2023;
		end
		32'h0000C78A: begin
				q			<=			16'h0007;
		end
		32'h0000C78C: begin
				q			<=			16'h8793;
		end
		32'h0000C78E: begin
				q			<=			16'hFFF7;
		end
		32'h0000C790: begin
				q			<=			16'hF06F;
		end
		32'h0000C792: begin
				q			<=			16'hFADF;
		end
		32'h0000C794: begin
				q			<=			16'h6A33;
		end
		32'h0000C796: begin
				q			<=			16'h016A;
		end
		32'h0000C798: begin
				q			<=			16'h6AB3;
		end
		32'h0000C79A: begin
				q			<=			16'h015A;
		end
		32'h0000C79C: begin
				q			<=			16'hEAB3;
		end
		32'h0000C79E: begin
				q			<=			16'h00FA;
		end
		32'h0000C7A0: begin
				q			<=			16'h0713;
		end
		32'h0000C7A2: begin
				q			<=			16'h0020;
		end
		32'h0000C7A4: begin
				q			<=			16'h8AE3;
		end
		32'h0000C7A6: begin
				q			<=			16'hD20A;
		end
		32'h0000C7A8: begin
				q			<=			16'h0713;
		end
		32'h0000C7AA: begin
				q			<=			16'h0030;
		end
		32'h0000C7AC: begin
				q			<=			16'hF06F;
		end
		32'h0000C7AE: begin
				q			<=			16'hD2DF;
		end
		32'h0000C7B0: begin
				q			<=			16'h0513;
		end
		32'h0000C7B2: begin
				q			<=			16'h0000;
		end
		32'h0000C7B4: begin
				q			<=			16'h0713;
		end
		32'h0000C7B6: begin
				q			<=			16'h0010;
		end
		32'h0000C7B8: begin
				q			<=			16'hF06F;
		end
		32'h0000C7BA: begin
				q			<=			16'hD21F;
		end
		32'h0000C7BC: begin
				q			<=			16'h2703;
		end
		32'h0000C7BE: begin
				q			<=			16'h0301;
		end
		32'h0000C7C0: begin
				q			<=			16'h2E03;
		end
		32'h0000C7C2: begin
				q			<=			16'h0401;
		end
		32'h0000C7C4: begin
				q			<=			16'h0537;
		end
		32'h0000C7C6: begin
				q			<=			16'h0001;
		end
		32'h0000C7C8: begin
				q			<=			16'h0693;
		end
		32'h0000C7CA: begin
				q			<=			16'hFFF5;
		end
		32'h0000C7CC: begin
				q			<=			16'h5F93;
		end
		32'h0000C7CE: begin
				q			<=			16'h0107;
		end
		32'h0000C7D0: begin
				q			<=			16'h5A93;
		end
		32'h0000C7D2: begin
				q			<=			16'h010E;
		end
		32'h0000C7D4: begin
				q			<=			16'h7733;
		end
		32'h0000C7D6: begin
				q			<=			16'h00D7;
		end
		32'h0000C7D8: begin
				q			<=			16'h7E33;
		end
		32'h0000C7DA: begin
				q			<=			16'h00DE;
		end
		32'h0000C7DC: begin
				q			<=			16'h87B3;
		end
		32'h0000C7DE: begin
				q			<=			16'h02EA;
		end
		32'h0000C7E0: begin
				q			<=			16'h0633;
		end
		32'h0000C7E2: begin
				q			<=			16'h03C7;
		end
		32'h0000C7E4: begin
				q			<=			16'h8833;
		end
		32'h0000C7E6: begin
				q			<=			16'h03CF;
		end
		32'h0000C7E8: begin
				q			<=			16'h85B3;
		end
		32'h0000C7EA: begin
				q			<=			16'h0107;
		end
		32'h0000C7EC: begin
				q			<=			16'h5793;
		end
		32'h0000C7EE: begin
				q			<=			16'h0106;
		end
		32'h0000C7F0: begin
				q			<=			16'h87B3;
		end
		32'h0000C7F2: begin
				q			<=			16'h00B7;
		end
		32'h0000C7F4: begin
				q			<=			16'h8B33;
		end
		32'h0000C7F6: begin
				q			<=			16'h035F;
		end
		32'h0000C7F8: begin
				q			<=			16'hF463;
		end
		32'h0000C7FA: begin
				q			<=			16'h0107;
		end
		32'h0000C7FC: begin
				q			<=			16'h0B33;
		end
		32'h0000C7FE: begin
				q			<=			16'h00AB;
		end
		32'h0000C800: begin
				q			<=			16'h2F03;
		end
		32'h0000C802: begin
				q			<=			16'h0441;
		end
		32'h0000C804: begin
				q			<=			16'hD293;
		end
		32'h0000C806: begin
				q			<=			16'h0107;
		end
		32'h0000C808: begin
				q			<=			16'hF7B3;
		end
		32'h0000C80A: begin
				q			<=			16'h00D7;
		end
		32'h0000C80C: begin
				q			<=			16'h7633;
		end
		32'h0000C80E: begin
				q			<=			16'h00D6;
		end
		32'h0000C810: begin
				q			<=			16'h9793;
		end
		32'h0000C812: begin
				q			<=			16'h0107;
		end
		32'h0000C814: begin
				q			<=			16'h87B3;
		end
		32'h0000C816: begin
				q			<=			16'h00C7;
		end
		32'h0000C818: begin
				q			<=			16'h5493;
		end
		32'h0000C81A: begin
				q			<=			16'h010F;
		end
		32'h0000C81C: begin
				q			<=			16'h7F33;
		end
		32'h0000C81E: begin
				q			<=			16'h00DF;
		end
		32'h0000C820: begin
				q			<=			16'h2223;
		end
		32'h0000C822: begin
				q			<=			16'h02F1;
		end
		32'h0000C824: begin
				q			<=			16'h2023;
		end
		32'h0000C826: begin
				q			<=			16'h06F1;
		end
		32'h0000C828: begin
				q			<=			16'h06B3;
		end
		32'h0000C82A: begin
				q			<=			16'h03E7;
		end
		32'h0000C82C: begin
				q			<=			16'h87B3;
		end
		32'h0000C82E: begin
				q			<=			16'h02E4;
		end
		32'h0000C830: begin
				q			<=			16'h8633;
		end
		32'h0000C832: begin
				q			<=			16'h03EF;
		end
		32'h0000C834: begin
				q			<=			16'h8533;
		end
		32'h0000C836: begin
				q			<=			16'h00C7;
		end
		32'h0000C838: begin
				q			<=			16'hD793;
		end
		32'h0000C83A: begin
				q			<=			16'h0106;
		end
		32'h0000C83C: begin
				q			<=			16'h87B3;
		end
		32'h0000C83E: begin
				q			<=			16'h00A7;
		end
		32'h0000C840: begin
				q			<=			16'h8A33;
		end
		32'h0000C842: begin
				q			<=			16'h029F;
		end
		32'h0000C844: begin
				q			<=			16'hF663;
		end
		32'h0000C846: begin
				q			<=			16'h00C7;
		end
		32'h0000C848: begin
				q			<=			16'h0637;
		end
		32'h0000C84A: begin
				q			<=			16'h0001;
		end
		32'h0000C84C: begin
				q			<=			16'h0A33;
		end
		32'h0000C84E: begin
				q			<=			16'h00CA;
		end
		32'h0000C850: begin
				q			<=			16'h0637;
		end
		32'h0000C852: begin
				q			<=			16'h0001;
		end
		32'h0000C854: begin
				q			<=			16'h0593;
		end
		32'h0000C856: begin
				q			<=			16'hFFF6;
		end
		32'h0000C858: begin
				q			<=			16'hF533;
		end
		32'h0000C85A: begin
				q			<=			16'h00B7;
		end
		32'h0000C85C: begin
				q			<=			16'hDD93;
		end
		32'h0000C85E: begin
				q			<=			16'h0107;
		end
		32'h0000C860: begin
				q			<=			16'h2783;
		end
		32'h0000C862: begin
				q			<=			16'h0341;
		end
		32'h0000C864: begin
				q			<=			16'hF6B3;
		end
		32'h0000C866: begin
				q			<=			16'h00B6;
		end
		32'h0000C868: begin
				q			<=			16'h1513;
		end
		32'h0000C86A: begin
				q			<=			16'h0105;
		end
		32'h0000C86C: begin
				q			<=			16'hD913;
		end
		32'h0000C86E: begin
				q			<=			16'h0107;
		end
		32'h0000C870: begin
				q			<=			16'hF5B3;
		end
		32'h0000C872: begin
				q			<=			16'h00B7;
		end
		32'h0000C874: begin
				q			<=			16'h0533;
		end
		32'h0000C876: begin
				q			<=			16'h00D5;
		end
		32'h0000C878: begin
				q			<=			16'h87B3;
		end
		32'h0000C87A: begin
				q			<=			16'h02BA;
		end
		32'h0000C87C: begin
				q			<=			16'h82B3;
		end
		32'h0000C87E: begin
				q			<=			16'h00A2;
		end
		32'h0000C880: begin
				q			<=			16'h06B3;
		end
		32'h0000C882: begin
				q			<=			16'h02BE;
		end
		32'h0000C884: begin
				q			<=			16'h0333;
		end
		32'h0000C886: begin
				q			<=			16'h03C9;
		end
		32'h0000C888: begin
				q			<=			16'h8833;
		end
		32'h0000C88A: begin
				q			<=			16'h0067;
		end
		32'h0000C88C: begin
				q			<=			16'hD793;
		end
		32'h0000C88E: begin
				q			<=			16'h0106;
		end
		32'h0000C890: begin
				q			<=			16'h87B3;
		end
		32'h0000C892: begin
				q			<=			16'h0107;
		end
		32'h0000C894: begin
				q			<=			16'h88B3;
		end
		32'h0000C896: begin
				q			<=			16'h032A;
		end
		32'h0000C898: begin
				q			<=			16'hF463;
		end
		32'h0000C89A: begin
				q			<=			16'h0067;
		end
		32'h0000C89C: begin
				q			<=			16'h88B3;
		end
		32'h0000C89E: begin
				q			<=			16'h00C8;
		end
		32'h0000C8A0: begin
				q			<=			16'hD993;
		end
		32'h0000C8A2: begin
				q			<=			16'h0107;
		end
		32'h0000C8A4: begin
				q			<=			16'h89B3;
		end
		32'h0000C8A6: begin
				q			<=			16'h0119;
		end
		32'h0000C8A8: begin
				q			<=			16'h08B7;
		end
		32'h0000C8AA: begin
				q			<=			16'h0001;
		end
		32'h0000C8AC: begin
				q			<=			16'h8613;
		end
		32'h0000C8AE: begin
				q			<=			16'hFFF8;
		end
		32'h0000C8B0: begin
				q			<=			16'hF833;
		end
		32'h0000C8B2: begin
				q			<=			16'h00C7;
		end
		32'h0000C8B4: begin
				q			<=			16'hF6B3;
		end
		32'h0000C8B6: begin
				q			<=			16'h00C6;
		end
		32'h0000C8B8: begin
				q			<=			16'h1813;
		end
		32'h0000C8BA: begin
				q			<=			16'h0108;
		end
		32'h0000C8BC: begin
				q			<=			16'h0833;
		end
		32'h0000C8BE: begin
				q			<=			16'h00D8;
		end
		32'h0000C8C0: begin
				q			<=			16'h0633;
		end
		32'h0000C8C2: begin
				q			<=			16'h02BF;
		end
		32'h0000C8C4: begin
				q			<=			16'h07B3;
		end
		32'h0000C8C6: begin
				q			<=			16'h03E9;
		end
		32'h0000C8C8: begin
				q			<=			16'h5E93;
		end
		32'h0000C8CA: begin
				q			<=			16'h0106;
		end
		32'h0000C8CC: begin
				q			<=			16'h86B3;
		end
		32'h0000C8CE: begin
				q			<=			16'h02B4;
		end
		32'h0000C8D0: begin
				q			<=			16'h86B3;
		end
		32'h0000C8D2: begin
				q			<=			16'h00F6;
		end
		32'h0000C8D4: begin
				q			<=			16'h86B3;
		end
		32'h0000C8D6: begin
				q			<=			16'h00DE;
		end
		32'h0000C8D8: begin
				q			<=			16'h8333;
		end
		32'h0000C8DA: begin
				q			<=			16'h0324;
		end
		32'h0000C8DC: begin
				q			<=			16'hF463;
		end
		32'h0000C8DE: begin
				q			<=			16'h00F6;
		end
		32'h0000C8E0: begin
				q			<=			16'h0333;
		end
		32'h0000C8E2: begin
				q			<=			16'h0113;
		end
		32'h0000C8E4: begin
				q			<=			16'hD793;
		end
		32'h0000C8E6: begin
				q			<=			16'h0106;
		end
		32'h0000C8E8: begin
				q			<=			16'h2E83;
		end
		32'h0000C8EA: begin
				q			<=			16'h0481;
		end
		32'h0000C8EC: begin
				q			<=			16'h87B3;
		end
		32'h0000C8EE: begin
				q			<=			16'h0067;
		end
		32'h0000C8F0: begin
				q			<=			16'h03B7;
		end
		32'h0000C8F2: begin
				q			<=			16'h0001;
		end
		32'h0000C8F4: begin
				q			<=			16'h2423;
		end
		32'h0000C8F6: begin
				q			<=			16'h02F1;
		end
		32'h0000C8F8: begin
				q			<=			16'h8793;
		end
		32'h0000C8FA: begin
				q			<=			16'hFFF3;
		end
		32'h0000C8FC: begin
				q			<=			16'hD413;
		end
		32'h0000C8FE: begin
				q			<=			16'h010E;
		end
		32'h0000C900: begin
				q			<=			16'hFEB3;
		end
		32'h0000C902: begin
				q			<=			16'h00FE;
		end
		32'h0000C904: begin
				q			<=			16'h08B3;
		end
		32'h0000C906: begin
				q			<=			16'h02E4;
		end
		32'h0000C908: begin
				q			<=			16'h7633;
		end
		32'h0000C90A: begin
				q			<=			16'h00F6;
		end
		32'h0000C90C: begin
				q			<=			16'hF6B3;
		end
		32'h0000C90E: begin
				q			<=			16'h00F6;
		end
		32'h0000C910: begin
				q			<=			16'h9693;
		end
		32'h0000C912: begin
				q			<=			16'h0106;
		end
		32'h0000C914: begin
				q			<=			16'h86B3;
		end
		32'h0000C916: begin
				q			<=			16'h00C6;
		end
		32'h0000C918: begin
				q			<=			16'h0333;
		end
		32'h0000C91A: begin
				q			<=			16'h03D7;
		end
		32'h0000C91C: begin
				q			<=			16'h8BB3;
		end
		32'h0000C91E: begin
				q			<=			16'h03DF;
		end
		32'h0000C920: begin
				q			<=			16'h87B3;
		end
		32'h0000C922: begin
				q			<=			16'h0178;
		end
		32'h0000C924: begin
				q			<=			16'h5893;
		end
		32'h0000C926: begin
				q			<=			16'h0103;
		end
		32'h0000C928: begin
				q			<=			16'h88B3;
		end
		32'h0000C92A: begin
				q			<=			16'h00F8;
		end
		32'h0000C92C: begin
				q			<=			16'h8633;
		end
		32'h0000C92E: begin
				q			<=			16'h028F;
		end
		32'h0000C930: begin
				q			<=			16'hF463;
		end
		32'h0000C932: begin
				q			<=			16'h0178;
		end
		32'h0000C934: begin
				q			<=			16'h0633;
		end
		32'h0000C936: begin
				q			<=			16'h0076;
		end
		32'h0000C938: begin
				q			<=			16'hD793;
		end
		32'h0000C93A: begin
				q			<=			16'h0108;
		end
		32'h0000C93C: begin
				q			<=			16'h0C37;
		end
		32'h0000C93E: begin
				q			<=			16'h0001;
		end
		32'h0000C940: begin
				q			<=			16'h87B3;
		end
		32'h0000C942: begin
				q			<=			16'h00C7;
		end
		32'h0000C944: begin
				q			<=			16'h0613;
		end
		32'h0000C946: begin
				q			<=			16'hFFFC;
		end
		32'h0000C948: begin
				q			<=			16'h2623;
		end
		32'h0000C94A: begin
				q			<=			16'h02F1;
		end
		32'h0000C94C: begin
				q			<=			16'hF7B3;
		end
		32'h0000C94E: begin
				q			<=			16'h00C8;
		end
		32'h0000C950: begin
				q			<=			16'h2883;
		end
		32'h0000C952: begin
				q			<=			16'h0381;
		end
		32'h0000C954: begin
				q			<=			16'h7333;
		end
		32'h0000C956: begin
				q			<=			16'h00C3;
		end
		32'h0000C958: begin
				q			<=			16'h9793;
		end
		32'h0000C95A: begin
				q			<=			16'h0107;
		end
		32'h0000C95C: begin
				q			<=			16'hD393;
		end
		32'h0000C95E: begin
				q			<=			16'h0108;
		end
		32'h0000C960: begin
				q			<=			16'hF633;
		end
		32'h0000C962: begin
				q			<=			16'h00C8;
		end
		32'h0000C964: begin
				q			<=			16'h87B3;
		end
		32'h0000C966: begin
				q			<=			16'h0067;
		end
		32'h0000C968: begin
				q			<=			16'h08B3;
		end
		32'h0000C96A: begin
				q			<=			16'h02CE;
		end
		32'h0000C96C: begin
				q			<=			16'h8CB3;
		end
		32'h0000C96E: begin
				q			<=			16'h03C3;
		end
		32'h0000C970: begin
				q			<=			16'hDD13;
		end
		32'h0000C972: begin
				q			<=			16'h0108;
		end
		32'h0000C974: begin
				q			<=			16'h8333;
		end
		32'h0000C976: begin
				q			<=			16'h02CA;
		end
		32'h0000C978: begin
				q			<=			16'h0333;
		end
		32'h0000C97A: begin
				q			<=			16'h0193;
		end
		32'h0000C97C: begin
				q			<=			16'h0333;
		end
		32'h0000C97E: begin
				q			<=			16'h006D;
		end
		32'h0000C980: begin
				q			<=			16'h8BB3;
		end
		32'h0000C982: begin
				q			<=			16'h027A;
		end
		32'h0000C984: begin
				q			<=			16'h7463;
		end
		32'h0000C986: begin
				q			<=			16'h0193;
		end
		32'h0000C988: begin
				q			<=			16'h8BB3;
		end
		32'h0000C98A: begin
				q			<=			16'h018B;
		end
		32'h0000C98C: begin
				q			<=			16'h5C13;
		end
		32'h0000C98E: begin
				q			<=			16'h0103;
		end
		32'h0000C990: begin
				q			<=			16'h0BB3;
		end
		32'h0000C992: begin
				q			<=			16'h017C;
		end
		32'h0000C994: begin
				q			<=			16'h0C37;
		end
		32'h0000C996: begin
				q			<=			16'h0001;
		end
		32'h0000C998: begin
				q			<=			16'h02B3;
		end
		32'h0000C99A: begin
				q			<=			16'h005B;
		end
		32'h0000C99C: begin
				q			<=			16'h0C93;
		end
		32'h0000C99E: begin
				q			<=			16'hFFFC;
		end
		32'h0000C9A0: begin
				q			<=			16'hB533;
		end
		32'h0000C9A2: begin
				q			<=			16'h00A2;
		end
		32'h0000C9A4: begin
				q			<=			16'h7333;
		end
		32'h0000C9A6: begin
				q			<=			16'h0193;
		end
		32'h0000C9A8: begin
				q			<=			16'h8DB3;
		end
		32'h0000C9AA: begin
				q			<=			16'h00AD;
		end
		32'h0000C9AC: begin
				q			<=			16'h1313;
		end
		32'h0000C9AE: begin
				q			<=			16'h0103;
		end
		32'h0000C9B0: begin
				q			<=			16'hF8B3;
		end
		32'h0000C9B2: begin
				q			<=			16'h0198;
		end
		32'h0000C9B4: begin
				q			<=			16'h8A33;
		end
		32'h0000C9B6: begin
				q			<=			16'h014D;
		end
		32'h0000C9B8: begin
				q			<=			16'h08B3;
		end
		32'h0000C9BA: begin
				q			<=			16'h0113;
		end
		32'h0000C9BC: begin
				q			<=			16'h8333;
		end
		32'h0000C9BE: begin
				q			<=			16'h0102;
		end
		32'h0000C9C0: begin
				q			<=			16'h3833;
		end
		32'h0000C9C2: begin
				q			<=			16'h0103;
		end
		32'h0000C9C4: begin
				q			<=			16'h2A23;
		end
		32'h0000C9C6: begin
				q			<=			16'h0061;
		end
		32'h0000C9C8: begin
				q			<=			16'h2223;
		end
		32'h0000C9CA: begin
				q			<=			16'h0661;
		end
		32'h0000C9CC: begin
				q			<=			16'h0333;
		end
		32'h0000C9CE: begin
				q			<=			16'h013A;
		end
		32'h0000C9D0: begin
				q			<=			16'h0B33;
		end
		32'h0000C9D2: begin
				q			<=			16'h0103;
		end
		32'h0000C9D4: begin
				q			<=			16'h39B3;
		end
		32'h0000C9D6: begin
				q			<=			16'h0133;
		end
		32'h0000C9D8: begin
				q			<=			16'h3833;
		end
		32'h0000C9DA: begin
				q			<=			16'h010B;
		end
		32'h0000C9DC: begin
				q			<=			16'hE833;
		end
		32'h0000C9DE: begin
				q			<=			16'h0109;
		end
		32'h0000C9E0: begin
				q			<=			16'h3533;
		end
		32'h0000C9E2: begin
				q			<=			16'h00AA;
		end
		32'h0000C9E4: begin
				q			<=			16'h0533;
		end
		32'h0000C9E6: begin
				q			<=			16'h00A8;
		end
		32'h0000C9E8: begin
				q			<=			16'h2803;
		end
		32'h0000C9EA: begin
				q			<=			16'h0281;
		end
		32'h0000C9EC: begin
				q			<=			16'h02B3;
		end
		32'h0000C9EE: begin
				q			<=			16'h00DB;
		end
		32'h0000C9F0: begin
				q			<=			16'h2983;
		end
		32'h0000C9F2: begin
				q			<=			16'h0281;
		end
		32'h0000C9F4: begin
				q			<=			16'hB6B3;
		end
		32'h0000C9F6: begin
				q			<=			16'h00D2;
		end
		32'h0000C9F8: begin
				q			<=			16'h0533;
		end
		32'h0000C9FA: begin
				q			<=			16'h0105;
		end
		32'h0000C9FC: begin
				q			<=			16'h2303;
		end
		32'h0000C9FE: begin
				q			<=			16'h02C1;
		end
		32'h0000CA00: begin
				q			<=			16'h0833;
		end
		32'h0000CA02: begin
				q			<=			16'h00D5;
		end
		32'h0000CA04: begin
				q			<=			16'h82B3;
		end
		32'h0000CA06: begin
				q			<=			16'h00F2;
		end
		32'h0000CA08: begin
				q			<=			16'h3533;
		end
		32'h0000CA0A: begin
				q			<=			16'h0135;
		end
		32'h0000CA0C: begin
				q			<=			16'h36B3;
		end
		32'h0000CA0E: begin
				q			<=			16'h00D8;
		end
		32'h0000CA10: begin
				q			<=			16'hB7B3;
		end
		32'h0000CA12: begin
				q			<=			16'h00F2;
		end
		32'h0000CA14: begin
				q			<=			16'h0DB3;
		end
		32'h0000CA16: begin
				q			<=			16'h0068;
		end
		32'h0000CA18: begin
				q			<=			16'h66B3;
		end
		32'h0000CA1A: begin
				q			<=			16'h00D5;
		end
		32'h0000CA1C: begin
				q			<=			16'h2503;
		end
		32'h0000CA1E: begin
				q			<=			16'h02C1;
		end
		32'h0000CA20: begin
				q			<=			16'h8333;
		end
		32'h0000CA22: begin
				q			<=			16'h00FD;
		end
		32'h0000CA24: begin
				q			<=			16'h82B3;
		end
		32'h0000CA26: begin
				q			<=			16'h0112;
		end
		32'h0000CA28: begin
				q			<=			16'hB8B3;
		end
		32'h0000CA2A: begin
				q			<=			16'h0112;
		end
		32'h0000CA2C: begin
				q			<=			16'h37B3;
		end
		32'h0000CA2E: begin
				q			<=			16'h00F3;
		end
		32'h0000CA30: begin
				q			<=			16'h2C23;
		end
		32'h0000CA32: begin
				q			<=			16'h0051;
		end
		32'h0000CA34: begin
				q			<=			16'h2423;
		end
		32'h0000CA36: begin
				q			<=			16'h0651;
		end
		32'h0000CA38: begin
				q			<=			16'h02B3;
		end
		32'h0000CA3A: begin
				q			<=			16'h0173;
		end
		32'h0000CA3C: begin
				q			<=			16'h2303;
		end
		32'h0000CA3E: begin
				q			<=			16'h04C1;
		end
		32'h0000CA40: begin
				q			<=			16'h8D33;
		end
		32'h0000CA42: begin
				q			<=			16'h0112;
		end
		32'h0000CA44: begin
				q			<=			16'hBDB3;
		end
		32'h0000CA46: begin
				q			<=			16'h00AD;
		end
		32'h0000CA48: begin
				q			<=			16'hE7B3;
		end
		32'h0000CA4A: begin
				q			<=			16'h00FD;
		end
		32'h0000CA4C: begin
				q			<=			16'hBBB3;
		end
		32'h0000CA4E: begin
				q			<=			16'h0172;
		end
		32'h0000CA50: begin
				q			<=			16'h38B3;
		end
		32'h0000CA52: begin
				q			<=			16'h011D;
		end
		32'h0000CA54: begin
				q			<=			16'h86B3;
		end
		32'h0000CA56: begin
				q			<=			16'h00F6;
		end
		32'h0000CA58: begin
				q			<=			16'h5293;
		end
		32'h0000CA5A: begin
				q			<=			16'h0103;
		end
		32'h0000CA5C: begin
				q			<=			16'hEA33;
		end
		32'h0000CA5E: begin
				q			<=			16'h011B;
		end
		32'h0000CA60: begin
				q			<=			16'h7333;
		end
		32'h0000CA62: begin
				q			<=			16'h0193;
		end
		32'h0000CA64: begin
				q			<=			16'h07B3;
		end
		32'h0000CA66: begin
				q			<=			16'h0267;
		end
		32'h0000CA68: begin
				q			<=			16'h8A33;
		end
		32'h0000CA6A: begin
				q			<=			16'h0146;
		end
		32'h0000CA6C: begin
				q			<=			16'h8733;
		end
		32'h0000CA6E: begin
				q			<=			16'h02E2;
		end
		32'h0000CA70: begin
				q			<=			16'hD893;
		end
		32'h0000CA72: begin
				q			<=			16'h0107;
		end
		32'h0000CA74: begin
				q			<=			16'h86B3;
		end
		32'h0000CA76: begin
				q			<=			16'h026F;
		end
		32'h0000CA78: begin
				q			<=			16'h0733;
		end
		32'h0000CA7A: begin
				q			<=			16'h00D7;
		end
		32'h0000CA7C: begin
				q			<=			16'h88B3;
		end
		32'h0000CA7E: begin
				q			<=			16'h00E8;
		end
		32'h0000CA80: begin
				q			<=			16'h8FB3;
		end
		32'h0000CA82: begin
				q			<=			16'h025F;
		end
		32'h0000CA84: begin
				q			<=			16'hF463;
		end
		32'h0000CA86: begin
				q			<=			16'h00D8;
		end
		32'h0000CA88: begin
				q			<=			16'h8FB3;
		end
		32'h0000CA8A: begin
				q			<=			16'h018F;
		end
		32'h0000CA8C: begin
				q			<=			16'h2983;
		end
		32'h0000CA8E: begin
				q			<=			16'h03C1;
		end
		32'h0000CA90: begin
				q			<=			16'h06B7;
		end
		32'h0000CA92: begin
				q			<=			16'h0001;
		end
		32'h0000CA94: begin
				q			<=			16'h8513;
		end
		32'h0000CA96: begin
				q			<=			16'hFFF6;
		end
		32'h0000CA98: begin
				q			<=			16'hD713;
		end
		32'h0000CA9A: begin
				q			<=			16'h0108;
		end
		32'h0000CA9C: begin
				q			<=			16'hF8B3;
		end
		32'h0000CA9E: begin
				q			<=			16'h00A8;
		end
		32'h0000CAA0: begin
				q			<=			16'h0733;
		end
		32'h0000CAA2: begin
				q			<=			16'h01F7;
		end
		32'h0000CAA4: begin
				q			<=			16'hF7B3;
		end
		32'h0000CAA6: begin
				q			<=			16'h00A7;
		end
		32'h0000CAA8: begin
				q			<=			16'hDF93;
		end
		32'h0000CAAA: begin
				q			<=			16'h0109;
		end
		32'h0000CAAC: begin
				q			<=			16'h9893;
		end
		32'h0000CAAE: begin
				q			<=			16'h0108;
		end
		32'h0000CAB0: begin
				q			<=			16'hF9B3;
		end
		32'h0000CAB2: begin
				q			<=			16'h00A9;
		end
		32'h0000CAB4: begin
				q			<=			16'h88B3;
		end
		32'h0000CAB6: begin
				q			<=			16'h00F8;
		end
		32'h0000CAB8: begin
				q			<=			16'h8B33;
		end
		32'h0000CABA: begin
				q			<=			16'h03FA;
		end
		32'h0000CABC: begin
				q			<=			16'h0D93;
		end
		32'h0000CABE: begin
				q			<=			16'h0007;
		end
		32'h0000CAC0: begin
				q			<=			16'h07B3;
		end
		32'h0000CAC2: begin
				q			<=			16'h033E;
		end
		32'h0000CAC4: begin
				q			<=			16'h8AB3;
		end
		32'h0000CAC6: begin
				q			<=			16'h033A;
		end
		32'h0000CAC8: begin
				q			<=			16'hD813;
		end
		32'h0000CACA: begin
				q			<=			16'h0107;
		end
		32'h0000CACC: begin
				q			<=			16'h8E33;
		end
		32'h0000CACE: begin
				q			<=			16'h03CF;
		end
		32'h0000CAD0: begin
				q			<=			16'h8AB3;
		end
		32'h0000CAD2: begin
				q			<=			16'h01CA;
		end
		32'h0000CAD4: begin
				q			<=			16'h0AB3;
		end
		32'h0000CAD6: begin
				q			<=			16'h0158;
		end
		32'h0000CAD8: begin
				q			<=			16'hF463;
		end
		32'h0000CADA: begin
				q			<=			16'h01CA;
		end
		32'h0000CADC: begin
				q			<=			16'h0B33;
		end
		32'h0000CADE: begin
				q			<=			16'h00DB;
		end
		32'h0000CAE0: begin
				q			<=			16'hD813;
		end
		32'h0000CAE2: begin
				q			<=			16'h010A;
		end
		32'h0000CAE4: begin
				q			<=			16'h0733;
		end
		32'h0000CAE6: begin
				q			<=			16'h0168;
		end
		32'h0000CAE8: begin
				q			<=			16'h0B37;
		end
		32'h0000CAEA: begin
				q			<=			16'h0001;
		end
		32'h0000CAEC: begin
				q			<=			16'h2423;
		end
		32'h0000CAEE: begin
				q			<=			16'h02E1;
		end
		32'h0000CAF0: begin
				q			<=			16'h0713;
		end
		32'h0000CAF2: begin
				q			<=			16'hFFFB;
		end
		32'h0000CAF4: begin
				q			<=			16'hF833;
		end
		32'h0000CAF6: begin
				q			<=			16'h00EA;
		end
		32'h0000CAF8: begin
				q			<=			16'hF7B3;
		end
		32'h0000CAFA: begin
				q			<=			16'h00E7;
		end
		32'h0000CAFC: begin
				q			<=			16'h1813;
		end
		32'h0000CAFE: begin
				q			<=			16'h0108;
		end
		32'h0000CB00: begin
				q			<=			16'h0833;
		end
		32'h0000CB02: begin
				q			<=			16'h00F8;
		end
		32'h0000CB04: begin
				q			<=			16'h86B3;
		end
		32'h0000CB06: begin
				q			<=			16'h03D5;
		end
		32'h0000CB08: begin
				q			<=			16'h0E33;
		end
		32'h0000CB0A: begin
				q			<=			16'h03D9;
		end
		32'h0000CB0C: begin
				q			<=			16'hD513;
		end
		32'h0000CB0E: begin
				q			<=			16'h0106;
		end
		32'h0000CB10: begin
				q			<=			16'h07B3;
		end
		32'h0000CB12: begin
				q			<=			16'h02B4;
		end
		32'h0000CB14: begin
				q			<=			16'h87B3;
		end
		32'h0000CB16: begin
				q			<=			16'h01C7;
		end
		32'h0000CB18: begin
				q			<=			16'h07B3;
		end
		32'h0000CB1A: begin
				q			<=			16'h00F5;
		end
		32'h0000CB1C: begin
				q			<=			16'h0733;
		end
		32'h0000CB1E: begin
				q			<=			16'h0289;
		end
		32'h0000CB20: begin
				q			<=			16'hF463;
		end
		32'h0000CB22: begin
				q			<=			16'h01C7;
		end
		32'h0000CB24: begin
				q			<=			16'h0733;
		end
		32'h0000CB26: begin
				q			<=			16'h0167;
		end
		32'h0000CB28: begin
				q			<=			16'hD513;
		end
		32'h0000CB2A: begin
				q			<=			16'h0107;
		end
		32'h0000CB2C: begin
				q			<=			16'h0733;
		end
		32'h0000CB2E: begin
				q			<=			16'h00E5;
		end
		32'h0000CB30: begin
				q			<=			16'h0B37;
		end
		32'h0000CB32: begin
				q			<=			16'h0001;
		end
		32'h0000CB34: begin
				q			<=			16'h2623;
		end
		32'h0000CB36: begin
				q			<=			16'h02E1;
		end
		32'h0000CB38: begin
				q			<=			16'h0713;
		end
		32'h0000CB3A: begin
				q			<=			16'hFFFB;
		end
		32'h0000CB3C: begin
				q			<=			16'hF533;
		end
		32'h0000CB3E: begin
				q			<=			16'h00E7;
		end
		32'h0000CB40: begin
				q			<=			16'hF6B3;
		end
		32'h0000CB42: begin
				q			<=			16'h00E6;
		end
		32'h0000CB44: begin
				q			<=			16'h8E33;
		end
		32'h0000CB46: begin
				q			<=			16'h03E3;
		end
		32'h0000CB48: begin
				q			<=			16'h1513;
		end
		32'h0000CB4A: begin
				q			<=			16'h0105;
		end
		32'h0000CB4C: begin
				q			<=			16'h0533;
		end
		32'h0000CB4E: begin
				q			<=			16'h00D5;
		end
		32'h0000CB50: begin
				q			<=			16'h0733;
		end
		32'h0000CB52: begin
				q			<=			16'h02CF;
		end
		32'h0000CB54: begin
				q			<=			16'h87B3;
		end
		32'h0000CB56: begin
				q			<=			16'h02C4;
		end
		32'h0000CB58: begin
				q			<=			16'h5693;
		end
		32'h0000CB5A: begin
				q			<=			16'h0107;
		end
		32'h0000CB5C: begin
				q			<=			16'h87B3;
		end
		32'h0000CB5E: begin
				q			<=			16'h01C7;
		end
		32'h0000CB60: begin
				q			<=			16'h87B3;
		end
		32'h0000CB62: begin
				q			<=			16'h00F6;
		end
		32'h0000CB64: begin
				q			<=			16'h8AB3;
		end
		32'h0000CB66: begin
				q			<=			16'h0274;
		end
		32'h0000CB68: begin
				q			<=			16'hF463;
		end
		32'h0000CB6A: begin
				q			<=			16'h01C7;
		end
		32'h0000CB6C: begin
				q			<=			16'h8AB3;
		end
		32'h0000CB6E: begin
				q			<=			16'h016A;
		end
		32'h0000CB70: begin
				q			<=			16'h06B7;
		end
		32'h0000CB72: begin
				q			<=			16'h0001;
		end
		32'h0000CB74: begin
				q			<=			16'h8E13;
		end
		32'h0000CB76: begin
				q			<=			16'hFFF6;
		end
		32'h0000CB78: begin
				q			<=			16'hF6B3;
		end
		32'h0000CB7A: begin
				q			<=			16'h01C7;
		end
		32'h0000CB7C: begin
				q			<=			16'hDB93;
		end
		32'h0000CB7E: begin
				q			<=			16'h0107;
		end
		32'h0000CB80: begin
				q			<=			16'h07B3;
		end
		32'h0000CB82: begin
				q			<=			16'h011D;
		end
		32'h0000CB84: begin
				q			<=			16'h7733;
		end
		32'h0000CB86: begin
				q			<=			16'h01C7;
		end
		32'h0000CB88: begin
				q			<=			16'hB8B3;
		end
		32'h0000CB8A: begin
				q			<=			16'h0117;
		end
		32'h0000CB8C: begin
				q			<=			16'h0A33;
		end
		32'h0000CB8E: begin
				q			<=			16'h01BA;
		end
		32'h0000CB90: begin
				q			<=			16'h9693;
		end
		32'h0000CB92: begin
				q			<=			16'h0106;
		end
		32'h0000CB94: begin
				q			<=			16'h86B3;
		end
		32'h0000CB96: begin
				q			<=			16'h00E6;
		end
		32'h0000CB98: begin
				q			<=			16'h0D33;
		end
		32'h0000CB9A: begin
				q			<=			16'h011A;
		end
		32'h0000CB9C: begin
				q			<=			16'h2703;
		end
		32'h0000CB9E: begin
				q			<=			16'h0281;
		end
		32'h0000CBA0: begin
				q			<=			16'h38B3;
		end
		32'h0000CBA2: begin
				q			<=			16'h011D;
		end
		32'h0000CBA4: begin
				q			<=			16'h3A33;
		end
		32'h0000CBA6: begin
				q			<=			16'h01BA;
		end
		32'h0000CBA8: begin
				q			<=			16'h87B3;
		end
		32'h0000CBAA: begin
				q			<=			16'h0107;
		end
		32'h0000CBAC: begin
				q			<=			16'h6A33;
		end
		32'h0000CBAE: begin
				q			<=			16'h011A;
		end
		32'h0000CBB0: begin
				q			<=			16'h2883;
		end
		32'h0000CBB2: begin
				q			<=			16'h0281;
		end
		32'h0000CBB4: begin
				q			<=			16'hB833;
		end
		32'h0000CBB6: begin
				q			<=			16'h0107;
		end
		32'h0000CBB8: begin
				q			<=			16'h0B33;
		end
		32'h0000CBBA: begin
				q			<=			16'h00ED;
		end
		32'h0000CBBC: begin
				q			<=			16'h2703;
		end
		32'h0000CBBE: begin
				q			<=			16'h02C1;
		end
		32'h0000CBC0: begin
				q			<=			16'h0CB3;
		end
		32'h0000CBC2: begin
				q			<=			16'h010B;
		end
		32'h0000CBC4: begin
				q			<=			16'h87B3;
		end
		32'h0000CBC6: begin
				q			<=			16'h00A7;
		end
		32'h0000CBC8: begin
				q			<=			16'h3B33;
		end
		32'h0000CBCA: begin
				q			<=			16'h011B;
		end
		32'h0000CBCC: begin
				q			<=			16'hB833;
		end
		32'h0000CBCE: begin
				q			<=			16'h010C;
		end
		32'h0000CBD0: begin
				q			<=			16'hB533;
		end
		32'h0000CBD2: begin
				q			<=			16'h00A7;
		end
		32'h0000CBD4: begin
				q			<=			16'h8733;
		end
		32'h0000CBD6: begin
				q			<=			16'h00EC;
		end
		32'h0000CBD8: begin
				q			<=			16'h6B33;
		end
		32'h0000CBDA: begin
				q			<=			16'h010B;
		end
		32'h0000CBDC: begin
				q			<=			16'h2803;
		end
		32'h0000CBDE: begin
				q			<=			16'h02C1;
		end
		32'h0000CBE0: begin
				q			<=			16'h0C33;
		end
		32'h0000CBE2: begin
				q			<=			16'h00A7;
		end
		32'h0000CBE4: begin
				q			<=			16'h8BB3;
		end
		32'h0000CBE6: begin
				q			<=			16'h015B;
		end
		32'h0000CBE8: begin
				q			<=			16'h87B3;
		end
		32'h0000CBEA: begin
				q			<=			16'h00D7;
		end
		32'h0000CBEC: begin
				q			<=			16'hB6B3;
		end
		32'h0000CBEE: begin
				q			<=			16'h00D7;
		end
		32'h0000CBF0: begin
				q			<=			16'h0AB3;
		end
		32'h0000CBF2: begin
				q			<=			16'h017C;
		end
		32'h0000CBF4: begin
				q			<=			16'h8E33;
		end
		32'h0000CBF6: begin
				q			<=			16'h00DA;
		end
		32'h0000CBF8: begin
				q			<=			16'h3733;
		end
		32'h0000CBFA: begin
				q			<=			16'h0107;
		end
		32'h0000CBFC: begin
				q			<=			16'h3533;
		end
		32'h0000CBFE: begin
				q			<=			16'h00AC;
		end
		32'h0000CC00: begin
				q			<=			16'h6733;
		end
		32'h0000CC02: begin
				q			<=			16'h00A7;
		end
		32'h0000CC04: begin
				q			<=			16'h36B3;
		end
		32'h0000CC06: begin
				q			<=			16'h00DE;
		end
		32'h0000CC08: begin
				q			<=			16'h0A33;
		end
		32'h0000CC0A: begin
				q			<=			16'h016A;
		end
		32'h0000CC0C: begin
				q			<=			16'hBAB3;
		end
		32'h0000CC0E: begin
				q			<=			16'h017A;
		end
		32'h0000CC10: begin
				q			<=			16'h0A33;
		end
		32'h0000CC12: begin
				q			<=			16'h00EA;
		end
		32'h0000CC14: begin
				q			<=			16'hEAB3;
		end
		32'h0000CC16: begin
				q			<=			16'h00DA;
		end
		32'h0000CC18: begin
				q			<=			16'h06B3;
		end
		32'h0000CC1A: begin
				q			<=			16'h015A;
		end
		32'h0000CC1C: begin
				q			<=			16'h8833;
		end
		32'h0000CC1E: begin
				q			<=			16'h02CE;
		end
		32'h0000CC20: begin
				q			<=			16'h2623;
		end
		32'h0000CC22: begin
				q			<=			16'h06F1;
		end
		32'h0000CC24: begin
				q			<=			16'h8A33;
		end
		32'h0000CC26: begin
				q			<=			16'h03D3;
		end
		32'h0000CC28: begin
				q			<=			16'h5513;
		end
		32'h0000CC2A: begin
				q			<=			16'h0108;
		end
		32'h0000CC2C: begin
				q			<=			16'h0733;
		end
		32'h0000CC2E: begin
				q			<=			16'h02C4;
		end
		32'h0000CC30: begin
				q			<=			16'h0733;
		end
		32'h0000CC32: begin
				q			<=			16'h0147;
		end
		32'h0000CC34: begin
				q			<=			16'h0733;
		end
		32'h0000CC36: begin
				q			<=			16'h00E5;
		end
		32'h0000CC38: begin
				q			<=			16'h08B3;
		end
		32'h0000CC3A: begin
				q			<=			16'h0274;
		end
		32'h0000CC3C: begin
				q			<=			16'h7663;
		end
		32'h0000CC3E: begin
				q			<=			16'h0147;
		end
		32'h0000CC40: begin
				q			<=			16'h0537;
		end
		32'h0000CC42: begin
				q			<=			16'h0001;
		end
		32'h0000CC44: begin
				q			<=			16'h88B3;
		end
		32'h0000CC46: begin
				q			<=			16'h00A8;
		end
		32'h0000CC48: begin
				q			<=			16'h0A37;
		end
		32'h0000CC4A: begin
				q			<=			16'h0001;
		end
		32'h0000CC4C: begin
				q			<=			16'h5513;
		end
		32'h0000CC4E: begin
				q			<=			16'h0107;
		end
		32'h0000CC50: begin
				q			<=			16'h0A93;
		end
		32'h0000CC52: begin
				q			<=			16'hFFFA;
		end
		32'h0000CC54: begin
				q			<=			16'h08B3;
		end
		32'h0000CC56: begin
				q			<=			16'h0115;
		end
		32'h0000CC58: begin
				q			<=			16'h7533;
		end
		32'h0000CC5A: begin
				q			<=			16'h0157;
		end
		32'h0000CC5C: begin
				q			<=			16'h7833;
		end
		32'h0000CC5E: begin
				q			<=			16'h0158;
		end
		32'h0000CC60: begin
				q			<=			16'h1513;
		end
		32'h0000CC62: begin
				q			<=			16'h0105;
		end
		32'h0000CC64: begin
				q			<=			16'h0AB3;
		end
		32'h0000CC66: begin
				q			<=			16'h0269;
		end
		32'h0000CC68: begin
				q			<=			16'h0533;
		end
		32'h0000CC6A: begin
				q			<=			16'h0105;
		end
		32'h0000CC6C: begin
				q			<=			16'h8833;
		end
		32'h0000CC6E: begin
				q			<=			16'h0265;
		end
		32'h0000CC70: begin
				q			<=			16'h85B3;
		end
		32'h0000CC72: begin
				q			<=			16'h02B2;
		end
		32'h0000CC74: begin
				q			<=			16'h5713;
		end
		32'h0000CC76: begin
				q			<=			16'h0108;
		end
		32'h0000CC78: begin
				q			<=			16'h85B3;
		end
		32'h0000CC7A: begin
				q			<=			16'h0155;
		end
		32'h0000CC7C: begin
				q			<=			16'h0733;
		end
		32'h0000CC7E: begin
				q			<=			16'h00B7;
		end
		32'h0000CC80: begin
				q			<=			16'h0933;
		end
		32'h0000CC82: begin
				q			<=			16'h0259;
		end
		32'h0000CC84: begin
				q			<=			16'h7463;
		end
		32'h0000CC86: begin
				q			<=			16'h0157;
		end
		32'h0000CC88: begin
				q			<=			16'h0933;
		end
		32'h0000CC8A: begin
				q			<=			16'h0149;
		end
		32'h0000CC8C: begin
				q			<=			16'h0AB7;
		end
		32'h0000CC8E: begin
				q			<=			16'h0001;
		end
		32'h0000CC90: begin
				q			<=			16'h5593;
		end
		32'h0000CC92: begin
				q			<=			16'h0107;
		end
		32'h0000CC94: begin
				q			<=			16'h8A13;
		end
		32'h0000CC96: begin
				q			<=			16'hFFFA;
		end
		32'h0000CC98: begin
				q			<=			16'h7833;
		end
		32'h0000CC9A: begin
				q			<=			16'h0148;
		end
		32'h0000CC9C: begin
				q			<=			16'h8933;
		end
		32'h0000CC9E: begin
				q			<=			16'h0125;
		end
		32'h0000CCA0: begin
				q			<=			16'h75B3;
		end
		32'h0000CCA2: begin
				q			<=			16'h0147;
		end
		32'h0000CCA4: begin
				q			<=			16'h9593;
		end
		32'h0000CCA6: begin
				q			<=			16'h0105;
		end
		32'h0000CCA8: begin
				q			<=			16'h0733;
		end
		32'h0000CCAA: begin
				q			<=			16'h033F;
		end
		32'h0000CCAC: begin
				q			<=			16'h85B3;
		end
		32'h0000CCAE: begin
				q			<=			16'h0105;
		end
		32'h0000CCB0: begin
				q			<=			16'h8F33;
		end
		32'h0000CCB2: begin
				q			<=			16'h03EF;
		end
		32'h0000CCB4: begin
				q			<=			16'h5813;
		end
		32'h0000CCB6: begin
				q			<=			16'h0107;
		end
		32'h0000CCB8: begin
				q			<=			16'h8A33;
		end
		32'h0000CCBA: begin
				q			<=			16'h03F4;
		end
		32'h0000CCBC: begin
				q			<=			16'h84B3;
		end
		32'h0000CCBE: begin
				q			<=			16'h0334;
		end
		32'h0000CCC0: begin
				q			<=			16'h84B3;
		end
		32'h0000CCC2: begin
				q			<=			16'h01E4;
		end
		32'h0000CCC4: begin
				q			<=			16'h04B3;
		end
		32'h0000CCC6: begin
				q			<=			16'h0098;
		end
		32'h0000CCC8: begin
				q			<=			16'hF463;
		end
		32'h0000CCCA: begin
				q			<=			16'h01E4;
		end
		32'h0000CCCC: begin
				q			<=			16'h0A33;
		end
		32'h0000CCCE: begin
				q			<=			16'h015A;
		end
		32'h0000CCD0: begin
				q			<=			16'hDB13;
		end
		32'h0000CCD2: begin
				q			<=			16'h0104;
		end
		32'h0000CCD4: begin
				q			<=			16'h0B33;
		end
		32'h0000CCD6: begin
				q			<=			16'h014B;
		end
		32'h0000CCD8: begin
				q			<=			16'h0A37;
		end
		32'h0000CCDA: begin
				q			<=			16'h0001;
		end
		32'h0000CCDC: begin
				q			<=			16'h0F13;
		end
		32'h0000CCDE: begin
				q			<=			16'hFFFA;
		end
		32'h0000CCE0: begin
				q			<=			16'hF833;
		end
		32'h0000CCE2: begin
				q			<=			16'h01E4;
		end
		32'h0000CCE4: begin
				q			<=			16'h7733;
		end
		32'h0000CCE6: begin
				q			<=			16'h01E7;
		end
		32'h0000CCE8: begin
				q			<=			16'h84B3;
		end
		32'h0000CCEA: begin
				q			<=			16'h0263;
		end
		32'h0000CCEC: begin
				q			<=			16'h1813;
		end
		32'h0000CCEE: begin
				q			<=			16'h0108;
		end
		32'h0000CCF0: begin
				q			<=			16'h0833;
		end
		32'h0000CCF2: begin
				q			<=			16'h00E8;
		end
		32'h0000CCF4: begin
				q			<=			16'h0F33;
		end
		32'h0000CCF6: begin
				q			<=			16'h0266;
		end
		32'h0000CCF8: begin
				q			<=			16'h8633;
		end
		32'h0000CCFA: begin
				q			<=			16'h02C2;
		end
		32'h0000CCFC: begin
				q			<=			16'h5713;
		end
		32'h0000CCFE: begin
				q			<=			16'h010F;
		end
		32'h0000CD00: begin
				q			<=			16'h0633;
		end
		32'h0000CD02: begin
				q			<=			16'h0096;
		end
		32'h0000CD04: begin
				q			<=			16'h0633;
		end
		32'h0000CD06: begin
				q			<=			16'h00C7;
		end
		32'h0000CD08: begin
				q			<=			16'h83B3;
		end
		32'h0000CD0A: begin
				q			<=			16'h0253;
		end
		32'h0000CD0C: begin
				q			<=			16'h7463;
		end
		32'h0000CD0E: begin
				q			<=			16'h0096;
		end
		32'h0000CD10: begin
				q			<=			16'h83B3;
		end
		32'h0000CD12: begin
				q			<=			16'h0143;
		end
		32'h0000CD14: begin
				q			<=			16'h0A37;
		end
		32'h0000CD16: begin
				q			<=			16'h0001;
		end
		32'h0000CD18: begin
				q			<=			16'h5713;
		end
		32'h0000CD1A: begin
				q			<=			16'h0106;
		end
		32'h0000CD1C: begin
				q			<=			16'h0493;
		end
		32'h0000CD1E: begin
				q			<=			16'hFFFA;
		end
		32'h0000CD20: begin
				q			<=			16'h03B3;
		end
		32'h0000CD22: begin
				q			<=			16'h0077;
		end
		32'h0000CD24: begin
				q			<=			16'h7733;
		end
		32'h0000CD26: begin
				q			<=			16'h0096;
		end
		32'h0000CD28: begin
				q			<=			16'h7F33;
		end
		32'h0000CD2A: begin
				q			<=			16'h009F;
		end
		32'h0000CD2C: begin
				q			<=			16'h1713;
		end
		32'h0000CD2E: begin
				q			<=			16'h0107;
		end
		32'h0000CD30: begin
				q			<=			16'h0733;
		end
		32'h0000CD32: begin
				q			<=			16'h01E7;
		end
		32'h0000CD34: begin
				q			<=			16'h0633;
		end
		32'h0000CD36: begin
				q			<=			16'h0334;
		end
		32'h0000CD38: begin
				q			<=			16'h8F33;
		end
		32'h0000CD3A: begin
				q			<=			16'h033E;
		end
		32'h0000CD3C: begin
				q			<=			16'h8EB3;
		end
		32'h0000CD3E: begin
				q			<=			16'h03DF;
		end
		32'h0000CD40: begin
				q			<=			16'h5A93;
		end
		32'h0000CD42: begin
				q			<=			16'h010F;
		end
		32'h0000CD44: begin
				q			<=			16'h0633;
		end
		32'h0000CD46: begin
				q			<=			16'h01D6;
		end
		32'h0000CD48: begin
				q			<=			16'h8633;
		end
		32'h0000CD4A: begin
				q			<=			16'h00CA;
		end
		32'h0000CD4C: begin
				q			<=			16'h04B3;
		end
		32'h0000CD4E: begin
				q			<=			16'h03F4;
		end
		32'h0000CD50: begin
				q			<=			16'h7463;
		end
		32'h0000CD52: begin
				q			<=			16'h01D6;
		end
		32'h0000CD54: begin
				q			<=			16'h84B3;
		end
		32'h0000CD56: begin
				q			<=			16'h0144;
		end
		32'h0000CD58: begin
				q			<=			16'h5C13;
		end
		32'h0000CD5A: begin
				q			<=			16'h0106;
		end
		32'h0000CD5C: begin
				q			<=			16'h0CB7;
		end
		32'h0000CD5E: begin
				q			<=			16'h0001;
		end
		32'h0000CD60: begin
				q			<=			16'h0C33;
		end
		32'h0000CD62: begin
				q			<=			16'h009C;
		end
		32'h0000CD64: begin
				q			<=			16'h0E33;
		end
		32'h0000CD66: begin
				q			<=			16'h00AE;
		end
		32'h0000CD68: begin
				q			<=			16'h8493;
		end
		32'h0000CD6A: begin
				q			<=			16'hFFFC;
		end
		32'h0000CD6C: begin
				q			<=			16'h3533;
		end
		32'h0000CD6E: begin
				q			<=			16'h00AE;
		end
		32'h0000CD70: begin
				q			<=			16'h86B3;
		end
		32'h0000CD72: begin
				q			<=			16'h0116;
		end
		32'h0000CD74: begin
				q			<=			16'h7633;
		end
		32'h0000CD76: begin
				q			<=			16'h0096;
		end
		32'h0000CD78: begin
				q			<=			16'h8DB3;
		end
		32'h0000CD7A: begin
				q			<=			16'h00A6;
		end
		32'h0000CD7C: begin
				q			<=			16'h7F33;
		end
		32'h0000CD7E: begin
				q			<=			16'h009F;
		end
		32'h0000CD80: begin
				q			<=			16'h0E33;
		end
		32'h0000CD82: begin
				q			<=			16'h00BE;
		end
		32'h0000CD84: begin
				q			<=			16'h1613;
		end
		32'h0000CD86: begin
				q			<=			16'h0106;
		end
		32'h0000CD88: begin
				q			<=			16'h0633;
		end
		32'h0000CD8A: begin
				q			<=			16'h01E6;
		end
		32'h0000CD8C: begin
				q			<=			16'h35B3;
		end
		32'h0000CD8E: begin
				q			<=			16'h00BE;
		end
		32'h0000CD90: begin
				q			<=			16'h8F33;
		end
		32'h0000CD92: begin
				q			<=			16'h012D;
		end
		32'h0000CD94: begin
				q			<=			16'h0E33;
		end
		32'h0000CD96: begin
				q			<=			16'h010E;
		end
		32'h0000CD98: begin
				q			<=			16'h0D33;
		end
		32'h0000CD9A: begin
				q			<=			16'h00BF;
		end
		32'h0000CD9C: begin
				q			<=			16'h0EB3;
		end
		32'h0000CD9E: begin
				q			<=			16'h016D;
		end
		32'h0000CDA0: begin
				q			<=			16'h2823;
		end
		32'h0000CDA2: begin
				q			<=			16'h07C1;
		end
		32'h0000CDA4: begin
				q			<=			16'h3E33;
		end
		32'h0000CDA6: begin
				q			<=			16'h010E;
		end
		32'h0000CDA8: begin
				q			<=			16'h8A33;
		end
		32'h0000CDAA: begin
				q			<=			16'h01CE;
		end
		32'h0000CDAC: begin
				q			<=			16'hB6B3;
		end
		32'h0000CDAE: begin
				q			<=			16'h0116;
		end
		32'h0000CDB0: begin
				q			<=			16'h35B3;
		end
		32'h0000CDB2: begin
				q			<=			16'h00BD;
		end
		32'h0000CDB4: begin
				q			<=			16'hB533;
		end
		32'h0000CDB6: begin
				q			<=			16'h00AD;
		end
		32'h0000CDB8: begin
				q			<=			16'h3933;
		end
		32'h0000CDBA: begin
				q			<=			16'h012F;
		end
		32'h0000CDBC: begin
				q			<=			16'hE533;
		end
		32'h0000CDBE: begin
				q			<=			16'h00A6;
		end
		32'h0000CDC0: begin
				q			<=			16'h6933;
		end
		32'h0000CDC2: begin
				q			<=			16'h00B9;
		end
		32'h0000CDC4: begin
				q			<=			16'hBEB3;
		end
		32'h0000CDC6: begin
				q			<=			16'h016E;
		end
		32'h0000CDC8: begin
				q			<=			16'h3E33;
		end
		32'h0000CDCA: begin
				q			<=			16'h01CA;
		end
		32'h0000CDCC: begin
				q			<=			16'h0533;
		end
		32'h0000CDCE: begin
				q			<=			16'h0125;
		end
		32'h0000CDD0: begin
				q			<=			16'hEEB3;
		end
		32'h0000CDD2: begin
				q			<=			16'h01CE;
		end
		32'h0000CDD4: begin
				q			<=			16'h0833;
		end
		32'h0000CDD6: begin
				q			<=			16'h00EA;
		end
		32'h0000CDD8: begin
				q			<=			16'h0533;
		end
		32'h0000CDDA: begin
				q			<=			16'h01D5;
		end
		32'h0000CDDC: begin
				q			<=			16'h3733;
		end
		32'h0000CDDE: begin
				q			<=			16'h00E8;
		end
		32'h0000CDE0: begin
				q			<=			16'h0533;
		end
		32'h0000CDE2: begin
				q			<=			16'h0075;
		end
		32'h0000CDE4: begin
				q			<=			16'h06B3;
		end
		32'h0000CDE6: begin
				q			<=			16'h00E5;
		end
		32'h0000CDE8: begin
				q			<=			16'h33B3;
		end
		32'h0000CDEA: begin
				q			<=			16'h0075;
		end
		32'h0000CDEC: begin
				q			<=			16'h0533;
		end
		32'h0000CDEE: begin
				q			<=			16'h0333;
		end
		32'h0000CDF0: begin
				q			<=			16'h0833;
		end
		32'h0000CDF2: begin
				q			<=			16'h00C8;
		end
		32'h0000CDF4: begin
				q			<=			16'hB733;
		end
		32'h0000CDF6: begin
				q			<=			16'h00E6;
		end
		32'h0000CDF8: begin
				q			<=			16'h3633;
		end
		32'h0000CDFA: begin
				q			<=			16'h00C8;
		end
		32'h0000CDFC: begin
				q			<=			16'h86B3;
		end
		32'h0000CDFE: begin
				q			<=			16'h0186;
		end
		32'h0000CE00: begin
				q			<=			16'h85B3;
		end
		32'h0000CE02: begin
				q			<=			16'h00C6;
		end
		32'h0000CE04: begin
				q			<=			16'hBC33;
		end
		32'h0000CE06: begin
				q			<=			16'h0186;
		end
		32'h0000CE08: begin
				q			<=			16'hB633;
		end
		32'h0000CE0A: begin
				q			<=			16'h00C5;
		end
		32'h0000CE0C: begin
				q			<=			16'h2A23;
		end
		32'h0000CE0E: begin
				q			<=			16'h0701;
		end
		32'h0000CE10: begin
				q			<=			16'hE733;
		end
		32'h0000CE12: begin
				q			<=			16'h00E3;
		end
		32'h0000CE14: begin
				q			<=			16'h8333;
		end
		32'h0000CE16: begin
				q			<=			16'h026F;
		end
		32'h0000CE18: begin
				q			<=			16'h5693;
		end
		32'h0000CE1A: begin
				q			<=			16'h0105;
		end
		32'h0000CE1C: begin
				q			<=			16'h6633;
		end
		32'h0000CE1E: begin
				q			<=			16'h00CC;
		end
		32'h0000CE20: begin
				q			<=			16'h89B3;
		end
		32'h0000CE22: begin
				q			<=			16'h0332;
		end
		32'h0000CE24: begin
				q			<=			16'h89B3;
		end
		32'h0000CE26: begin
				q			<=			16'h0069;
		end
		32'h0000CE28: begin
				q			<=			16'h8FB3;
		end
		32'h0000CE2A: begin
				q			<=			16'h03F2;
		end
		32'h0000CE2C: begin
				q			<=			16'h82B3;
		end
		32'h0000CE2E: begin
				q			<=			16'h0136;
		end
		32'h0000CE30: begin
				q			<=			16'hF463;
		end
		32'h0000CE32: begin
				q			<=			16'h0062;
		end
		32'h0000CE34: begin
				q			<=			16'h8FB3;
		end
		32'h0000CE36: begin
				q			<=			16'h019F;
		end
		32'h0000CE38: begin
				q			<=			16'hF6B3;
		end
		32'h0000CE3A: begin
				q			<=			16'h0092;
		end
		32'h0000CE3C: begin
				q			<=			16'h9693;
		end
		32'h0000CE3E: begin
				q			<=			16'h0106;
		end
		32'h0000CE40: begin
				q			<=			16'h74B3;
		end
		32'h0000CE42: begin
				q			<=			16'h0095;
		end
		32'h0000CE44: begin
				q			<=			16'h84B3;
		end
		32'h0000CE46: begin
				q			<=			16'h0096;
		end
		32'h0000CE48: begin
				q			<=			16'hD293;
		end
		32'h0000CE4A: begin
				q			<=			16'h0102;
		end
		32'h0000CE4C: begin
				q			<=			16'h85B3;
		end
		32'h0000CE4E: begin
				q			<=			16'h0095;
		end
		32'h0000CE50: begin
				q			<=			16'h82B3;
		end
		32'h0000CE52: begin
				q			<=			16'h00E2;
		end
		32'h0000CE54: begin
				q			<=			16'h2683;
		end
		32'h0000CE56: begin
				q			<=			16'h0141;
		end
		32'h0000CE58: begin
				q			<=			16'h2703;
		end
		32'h0000CE5A: begin
				q			<=			16'h0241;
		end
		32'h0000CE5C: begin
				q			<=			16'h82B3;
		end
		32'h0000CE5E: begin
				q			<=			16'h00C2;
		end
		32'h0000CE60: begin
				q			<=			16'hB4B3;
		end
		32'h0000CE62: begin
				q			<=			16'h0095;
		end
		32'h0000CE64: begin
				q			<=			16'h82B3;
		end
		32'h0000CE66: begin
				q			<=			16'h0092;
		end
		32'h0000CE68: begin
				q			<=			16'h8FB3;
		end
		32'h0000CE6A: begin
				q			<=			16'h01F2;
		end
		32'h0000CE6C: begin
				q			<=			16'h62B3;
		end
		32'h0000CE6E: begin
				q			<=			16'h00D7;
		end
		32'h0000CE70: begin
				q			<=			16'h2703;
		end
		32'h0000CE72: begin
				q			<=			16'h0181;
		end
		32'h0000CE74: begin
				q			<=			16'h9793;
		end
		32'h0000CE76: begin
				q			<=			16'h00D7;
		end
		32'h0000CE78: begin
				q			<=			16'h2E23;
		end
		32'h0000CE7A: begin
				q			<=			16'h07F1;
		end
		32'h0000CE7C: begin
				q			<=			16'h62B3;
		end
		32'h0000CE7E: begin
				q			<=			16'h0057;
		end
		32'h0000CE80: begin
				q			<=			16'h2C23;
		end
		32'h0000CE82: begin
				q			<=			16'h06B1;
		end
		32'h0000CE84: begin
				q			<=			16'hE7B3;
		end
		32'h0000CE86: begin
				q			<=			16'h0057;
		end
		32'h0000CE88: begin
				q			<=			16'h0713;
		end
		32'h0000CE8A: begin
				q			<=			16'h0601;
		end
		32'h0000CE8C: begin
				q			<=			16'h0613;
		end
		32'h0000CE8E: begin
				q			<=			16'h0000;
		end
		32'h0000CE90: begin
				q			<=			16'h0513;
		end
		32'h0000CE92: begin
				q			<=			16'h0040;
		end
		32'h0000CE94: begin
				q			<=			16'h2683;
		end
		32'h0000CE96: begin
				q			<=			16'h00C7;
		end
		32'h0000CE98: begin
				q			<=			16'h2583;
		end
		32'h0000CE9A: begin
				q			<=			16'h0107;
		end
		32'h0000CE9C: begin
				q			<=			16'h0613;
		end
		32'h0000CE9E: begin
				q			<=			16'h0016;
		end
		32'h0000CEA0: begin
				q			<=			16'hD693;
		end
		32'h0000CEA2: begin
				q			<=			16'h0136;
		end
		32'h0000CEA4: begin
				q			<=			16'h9593;
		end
		32'h0000CEA6: begin
				q			<=			16'h00D5;
		end
		32'h0000CEA8: begin
				q			<=			16'hE6B3;
		end
		32'h0000CEAA: begin
				q			<=			16'h00B6;
		end
		32'h0000CEAC: begin
				q			<=			16'h2023;
		end
		32'h0000CEAE: begin
				q			<=			16'h00D7;
		end
		32'h0000CEB0: begin
				q			<=			16'h0713;
		end
		32'h0000CEB2: begin
				q			<=			16'h0047;
		end
		32'h0000CEB4: begin
				q			<=			16'h10E3;
		end
		32'h0000CEB6: begin
				q			<=			16'hFEA6;
		end
		32'h0000CEB8: begin
				q			<=			16'h2703;
		end
		32'h0000CEBA: begin
				q			<=			16'h0601;
		end
		32'h0000CEBC: begin
				q			<=			16'h2683;
		end
		32'h0000CEBE: begin
				q			<=			16'h0681;
		end
		32'h0000CEC0: begin
				q			<=			16'h37B3;
		end
		32'h0000CEC2: begin
				q			<=			16'h00F0;
		end
		32'h0000CEC4: begin
				q			<=			16'hE7B3;
		end
		32'h0000CEC6: begin
				q			<=			16'h00E7;
		end
		32'h0000CEC8: begin
				q			<=			16'h2C23;
		end
		32'h0000CECA: begin
				q			<=			16'h04D1;
		end
		32'h0000CECC: begin
				q			<=			16'h2703;
		end
		32'h0000CECE: begin
				q			<=			16'h06C1;
		end
		32'h0000CED0: begin
				q			<=			16'h2683;
		end
		32'h0000CED2: begin
				q			<=			16'h0641;
		end
		32'h0000CED4: begin
				q			<=			16'h2823;
		end
		32'h0000CED6: begin
				q			<=			16'h04F1;
		end
		32'h0000CED8: begin
				q			<=			16'h2E23;
		end
		32'h0000CEDA: begin
				q			<=			16'h04E1;
		end
		32'h0000CEDC: begin
				q			<=			16'h2A23;
		end
		32'h0000CEDE: begin
				q			<=			16'h04D1;
		end
		32'h0000CEE0: begin
				q			<=			16'h1693;
		end
		32'h0000CEE2: begin
				q			<=			16'h00B7;
		end
		32'h0000CEE4: begin
				q			<=			16'hD463;
		end
		32'h0000CEE6: begin
				q			<=			16'h2406;
		end
		32'h0000CEE8: begin
				q			<=			16'h9793;
		end
		32'h0000CEEA: begin
				q			<=			16'h01F7;
		end
		32'h0000CEEC: begin
				q			<=			16'h0713;
		end
		32'h0000CEEE: begin
				q			<=			16'h0501;
		end
		32'h0000CEF0: begin
				q			<=			16'h0613;
		end
		32'h0000CEF2: begin
				q			<=			16'h0000;
		end
		32'h0000CEF4: begin
				q			<=			16'h0513;
		end
		32'h0000CEF6: begin
				q			<=			16'h0030;
		end
		32'h0000CEF8: begin
				q			<=			16'h2683;
		end
		32'h0000CEFA: begin
				q			<=			16'h0007;
		end
		32'h0000CEFC: begin
				q			<=			16'h2583;
		end
		32'h0000CEFE: begin
				q			<=			16'h0047;
		end
		32'h0000CF00: begin
				q			<=			16'h0613;
		end
		32'h0000CF02: begin
				q			<=			16'h0016;
		end
		32'h0000CF04: begin
				q			<=			16'hD693;
		end
		32'h0000CF06: begin
				q			<=			16'h0016;
		end
		32'h0000CF08: begin
				q			<=			16'h9593;
		end
		32'h0000CF0A: begin
				q			<=			16'h01F5;
		end
		32'h0000CF0C: begin
				q			<=			16'hE6B3;
		end
		32'h0000CF0E: begin
				q			<=			16'h00B6;
		end
		32'h0000CF10: begin
				q			<=			16'h2023;
		end
		32'h0000CF12: begin
				q			<=			16'h00D7;
		end
		32'h0000CF14: begin
				q			<=			16'h0713;
		end
		32'h0000CF16: begin
				q			<=			16'h0047;
		end
		32'h0000CF18: begin
				q			<=			16'h10E3;
		end
		32'h0000CF1A: begin
				q			<=			16'hFEA6;
		end
		32'h0000CF1C: begin
				q			<=			16'h2703;
		end
		32'h0000CF1E: begin
				q			<=			16'h05C1;
		end
		32'h0000CF20: begin
				q			<=			16'h37B3;
		end
		32'h0000CF22: begin
				q			<=			16'h00F0;
		end
		32'h0000CF24: begin
				q			<=			16'h5713;
		end
		32'h0000CF26: begin
				q			<=			16'h0017;
		end
		32'h0000CF28: begin
				q			<=			16'h2E23;
		end
		32'h0000CF2A: begin
				q			<=			16'h04E1;
		end
		32'h0000CF2C: begin
				q			<=			16'h2703;
		end
		32'h0000CF2E: begin
				q			<=			16'h0501;
		end
		32'h0000CF30: begin
				q			<=			16'h67B3;
		end
		32'h0000CF32: begin
				q			<=			16'h00F7;
		end
		32'h0000CF34: begin
				q			<=			16'h2823;
		end
		32'h0000CF36: begin
				q			<=			16'h04F1;
		end
		32'h0000CF38: begin
				q			<=			16'h2703;
		end
		32'h0000CF3A: begin
				q			<=			16'h01C1;
		end
		32'h0000CF3C: begin
				q			<=			16'h47B7;
		end
		32'h0000CF3E: begin
				q			<=			16'h0000;
		end
		32'h0000CF40: begin
				q			<=			16'h8793;
		end
		32'h0000CF42: begin
				q			<=			16'hFFF7;
		end
		32'h0000CF44: begin
				q			<=			16'h07B3;
		end
		32'h0000CF46: begin
				q			<=			16'h00F7;
		end
		32'h0000CF48: begin
				q			<=			16'h5463;
		end
		32'h0000CF4A: begin
				q			<=			16'h20F0;
		end
		32'h0000CF4C: begin
				q			<=			16'h2703;
		end
		32'h0000CF4E: begin
				q			<=			16'h0501;
		end
		32'h0000CF50: begin
				q			<=			16'h7693;
		end
		32'h0000CF52: begin
				q			<=			16'h0077;
		end
		32'h0000CF54: begin
				q			<=			16'h8463;
		end
		32'h0000CF56: begin
				q			<=			16'h0406;
		end
		32'h0000CF58: begin
				q			<=			16'h7693;
		end
		32'h0000CF5A: begin
				q			<=			16'h00F7;
		end
		32'h0000CF5C: begin
				q			<=			16'h0613;
		end
		32'h0000CF5E: begin
				q			<=			16'h0040;
		end
		32'h0000CF60: begin
				q			<=			16'h8E63;
		end
		32'h0000CF62: begin
				q			<=			16'h02C6;
		end
		32'h0000CF64: begin
				q			<=			16'h2683;
		end
		32'h0000CF66: begin
				q			<=			16'h0541;
		end
		32'h0000CF68: begin
				q			<=			16'h0713;
		end
		32'h0000CF6A: begin
				q			<=			16'h0047;
		end
		32'h0000CF6C: begin
				q			<=			16'h2823;
		end
		32'h0000CF6E: begin
				q			<=			16'h04E1;
		end
		32'h0000CF70: begin
				q			<=			16'h3713;
		end
		32'h0000CF72: begin
				q			<=			16'h0047;
		end
		32'h0000CF74: begin
				q			<=			16'h06B3;
		end
		32'h0000CF76: begin
				q			<=			16'h00D7;
		end
		32'h0000CF78: begin
				q			<=			16'hB733;
		end
		32'h0000CF7A: begin
				q			<=			16'h00E6;
		end
		32'h0000CF7C: begin
				q			<=			16'h2A23;
		end
		32'h0000CF7E: begin
				q			<=			16'h04D1;
		end
		32'h0000CF80: begin
				q			<=			16'h2683;
		end
		32'h0000CF82: begin
				q			<=			16'h0581;
		end
		32'h0000CF84: begin
				q			<=			16'h06B3;
		end
		32'h0000CF86: begin
				q			<=			16'h00D7;
		end
		32'h0000CF88: begin
				q			<=			16'h2C23;
		end
		32'h0000CF8A: begin
				q			<=			16'h04D1;
		end
		32'h0000CF8C: begin
				q			<=			16'hB6B3;
		end
		32'h0000CF8E: begin
				q			<=			16'h00E6;
		end
		32'h0000CF90: begin
				q			<=			16'h2703;
		end
		32'h0000CF92: begin
				q			<=			16'h05C1;
		end
		32'h0000CF94: begin
				q			<=			16'h86B3;
		end
		32'h0000CF96: begin
				q			<=			16'h00E6;
		end
		32'h0000CF98: begin
				q			<=			16'h2E23;
		end
		32'h0000CF9A: begin
				q			<=			16'h04D1;
		end
		32'h0000CF9C: begin
				q			<=			16'h2703;
		end
		32'h0000CF9E: begin
				q			<=			16'h05C1;
		end
		32'h0000CFA0: begin
				q			<=			16'h1693;
		end
		32'h0000CFA2: begin
				q			<=			16'h00B7;
		end
		32'h0000CFA4: begin
				q			<=			16'hD063;
		end
		32'h0000CFA6: begin
				q			<=			16'h0206;
		end
		32'h0000CFA8: begin
				q			<=			16'h07B7;
		end
		32'h0000CFAA: begin
				q			<=			16'hFFF0;
		end
		32'h0000CFAC: begin
				q			<=			16'h8793;
		end
		32'h0000CFAE: begin
				q			<=			16'hFFF7;
		end
		32'h0000CFB0: begin
				q			<=			16'h7733;
		end
		32'h0000CFB2: begin
				q			<=			16'h00F7;
		end
		32'h0000CFB4: begin
				q			<=			16'h2E23;
		end
		32'h0000CFB6: begin
				q			<=			16'h04E1;
		end
		32'h0000CFB8: begin
				q			<=			16'h2703;
		end
		32'h0000CFBA: begin
				q			<=			16'h01C1;
		end
		32'h0000CFBC: begin
				q			<=			16'h47B7;
		end
		32'h0000CFBE: begin
				q			<=			16'h0000;
		end
		32'h0000CFC0: begin
				q			<=			16'h07B3;
		end
		32'h0000CFC2: begin
				q			<=			16'h00F7;
		end
		32'h0000CFC4: begin
				q			<=			16'h0713;
		end
		32'h0000CFC6: begin
				q			<=			16'h0501;
		end
		32'h0000CFC8: begin
				q			<=			16'h0613;
		end
		32'h0000CFCA: begin
				q			<=			16'h0000;
		end
		32'h0000CFCC: begin
				q			<=			16'h0513;
		end
		32'h0000CFCE: begin
				q			<=			16'h0030;
		end
		32'h0000CFD0: begin
				q			<=			16'h2683;
		end
		32'h0000CFD2: begin
				q			<=			16'h0007;
		end
		32'h0000CFD4: begin
				q			<=			16'h2583;
		end
		32'h0000CFD6: begin
				q			<=			16'h0047;
		end
		32'h0000CFD8: begin
				q			<=			16'h0613;
		end
		32'h0000CFDA: begin
				q			<=			16'h0016;
		end
		32'h0000CFDC: begin
				q			<=			16'hD693;
		end
		32'h0000CFDE: begin
				q			<=			16'h0036;
		end
		32'h0000CFE0: begin
				q			<=			16'h9593;
		end
		32'h0000CFE2: begin
				q			<=			16'h01D5;
		end
		32'h0000CFE4: begin
				q			<=			16'hE6B3;
		end
		32'h0000CFE6: begin
				q			<=			16'h00B6;
		end
		32'h0000CFE8: begin
				q			<=			16'h2023;
		end
		32'h0000CFEA: begin
				q			<=			16'h00D7;
		end
		32'h0000CFEC: begin
				q			<=			16'h0713;
		end
		32'h0000CFEE: begin
				q			<=			16'h0047;
		end
		32'h0000CFF0: begin
				q			<=			16'h10E3;
		end
		32'h0000CFF2: begin
				q			<=			16'hFEA6;
		end
		32'h0000CFF4: begin
				q			<=			16'h8737;
		end
		32'h0000CFF6: begin
				q			<=			16'h0000;
		end
		32'h0000CFF8: begin
				q			<=			16'h0693;
		end
		32'h0000CFFA: begin
				q			<=			16'hFFE7;
		end
		32'h0000CFFC: begin
				q			<=			16'hCE63;
		end
		32'h0000CFFE: begin
				q			<=			16'h12F6;
		end
		32'h0000D000: begin
				q			<=			16'h2703;
		end
		32'h0000D002: begin
				q			<=			16'h05C1;
		end
		32'h0000D004: begin
				q			<=			16'h5713;
		end
		32'h0000D006: begin
				q			<=			16'h0037;
		end
		32'h0000D008: begin
				q			<=			16'h2E23;
		end
		32'h0000D00A: begin
				q			<=			16'h04E1;
		end
		32'h0000D00C: begin
				q			<=			16'h2703;
		end
		32'h0000D00E: begin
				q			<=			16'h05C1;
		end
		32'h0000D010: begin
				q			<=			16'h86B7;
		end
		32'h0000D012: begin
				q			<=			16'hFFFF;
		end
		32'h0000D014: begin
				q			<=			16'h2083;
		end
		32'h0000D016: begin
				q			<=			16'h0BC1;
		end
		32'h0000D018: begin
				q			<=			16'h1623;
		end
		32'h0000D01A: begin
				q			<=			16'h06E1;
		end
		32'h0000D01C: begin
				q			<=			16'h8737;
		end
		32'h0000D01E: begin
				q			<=			16'h0000;
		end
		32'h0000D020: begin
				q			<=			16'h0713;
		end
		32'h0000D022: begin
				q			<=			16'hFFF7;
		end
		32'h0000D024: begin
				q			<=			16'hF7B3;
		end
		32'h0000D026: begin
				q			<=			16'h00E7;
		end
		32'h0000D028: begin
				q			<=			16'h5703;
		end
		32'h0000D02A: begin
				q			<=			16'h06E1;
		end
		32'h0000D02C: begin
				q			<=			16'h2403;
		end
		32'h0000D02E: begin
				q			<=			16'h0B81;
		end
		32'h0000D030: begin
				q			<=			16'h2483;
		end
		32'h0000D032: begin
				q			<=			16'h0B41;
		end
		32'h0000D034: begin
				q			<=			16'h7733;
		end
		32'h0000D036: begin
				q			<=			16'h00D7;
		end
		32'h0000D038: begin
				q			<=			16'h67B3;
		end
		32'h0000D03A: begin
				q			<=			16'h00F7;
		end
		32'h0000D03C: begin
				q			<=			16'h1723;
		end
		32'h0000D03E: begin
				q			<=			16'h06F1;
		end
		32'h0000D040: begin
				q			<=			16'hD713;
		end
		32'h0000D042: begin
				q			<=			16'h0087;
		end
		32'h0000D044: begin
				q			<=			16'h2783;
		end
		32'h0000D046: begin
				q			<=			16'h0101;
		end
		32'h0000D048: begin
				q			<=			16'h7713;
		end
		32'h0000D04A: begin
				q			<=			16'h07F7;
		end
		32'h0000D04C: begin
				q			<=			16'h2903;
		end
		32'h0000D04E: begin
				q			<=			16'h0B01;
		end
		32'h0000D050: begin
				q			<=			16'h9793;
		end
		32'h0000D052: begin
				q			<=			16'h0077;
		end
		32'h0000D054: begin
				q			<=			16'h67B3;
		end
		32'h0000D056: begin
				q			<=			16'h00F7;
		end
		32'h0000D058: begin
				q			<=			16'h07A3;
		end
		32'h0000D05A: begin
				q			<=			16'h06F1;
		end
		32'h0000D05C: begin
				q			<=			16'h2703;
		end
		32'h0000D05E: begin
				q			<=			16'h00C1;
		end
		32'h0000D060: begin
				q			<=			16'h2783;
		end
		32'h0000D062: begin
				q			<=			16'h0501;
		end
		32'h0000D064: begin
				q			<=			16'h2983;
		end
		32'h0000D066: begin
				q			<=			16'h0AC1;
		end
		32'h0000D068: begin
				q			<=			16'h2A03;
		end
		32'h0000D06A: begin
				q			<=			16'h0A81;
		end
		32'h0000D06C: begin
				q			<=			16'h2023;
		end
		32'h0000D06E: begin
				q			<=			16'h00F7;
		end
		32'h0000D070: begin
				q			<=			16'h2783;
		end
		32'h0000D072: begin
				q			<=			16'h0541;
		end
		32'h0000D074: begin
				q			<=			16'h2A83;
		end
		32'h0000D076: begin
				q			<=			16'h0A41;
		end
		32'h0000D078: begin
				q			<=			16'h2B03;
		end
		32'h0000D07A: begin
				q			<=			16'h0A01;
		end
		32'h0000D07C: begin
				q			<=			16'h2223;
		end
		32'h0000D07E: begin
				q			<=			16'h00F7;
		end
		32'h0000D080: begin
				q			<=			16'h2783;
		end
		32'h0000D082: begin
				q			<=			16'h0581;
		end
		32'h0000D084: begin
				q			<=			16'h2B83;
		end
		32'h0000D086: begin
				q			<=			16'h09C1;
		end
		32'h0000D088: begin
				q			<=			16'h2C03;
		end
		32'h0000D08A: begin
				q			<=			16'h0981;
		end
		32'h0000D08C: begin
				q			<=			16'h2423;
		end
		32'h0000D08E: begin
				q			<=			16'h00F7;
		end
		32'h0000D090: begin
				q			<=			16'h2783;
		end
		32'h0000D092: begin
				q			<=			16'h06C1;
		end
		32'h0000D094: begin
				q			<=			16'h2C83;
		end
		32'h0000D096: begin
				q			<=			16'h0941;
		end
		32'h0000D098: begin
				q			<=			16'h2D03;
		end
		32'h0000D09A: begin
				q			<=			16'h0901;
		end
		32'h0000D09C: begin
				q			<=			16'h2623;
		end
		32'h0000D09E: begin
				q			<=			16'h00F7;
		end
		32'h0000D0A0: begin
				q			<=			16'h2D83;
		end
		32'h0000D0A2: begin
				q			<=			16'h08C1;
		end
		32'h0000D0A4: begin
				q			<=			16'h0513;
		end
		32'h0000D0A6: begin
				q			<=			16'h0007;
		end
		32'h0000D0A8: begin
				q			<=			16'h0113;
		end
		32'h0000D0AA: begin
				q			<=			16'h0C01;
		end
		32'h0000D0AC: begin
				q			<=			16'h8067;
		end
		32'h0000D0AE: begin
				q			<=			16'h0000;
		end
		32'h0000D0B0: begin
				q			<=			16'h2823;
		end
		32'h0000D0B2: begin
				q			<=			16'h0131;
		end
		32'h0000D0B4: begin
				q			<=			16'h2783;
		end
		32'h0000D0B6: begin
				q			<=			16'h0301;
		end
		32'h0000D0B8: begin
				q			<=			16'h2823;
		end
		32'h0000D0BA: begin
				q			<=			16'h04F1;
		end
		32'h0000D0BC: begin
				q			<=			16'h2783;
		end
		32'h0000D0BE: begin
				q			<=			16'h0341;
		end
		32'h0000D0C0: begin
				q			<=			16'h2A23;
		end
		32'h0000D0C2: begin
				q			<=			16'h04F1;
		end
		32'h0000D0C4: begin
				q			<=			16'h2783;
		end
		32'h0000D0C6: begin
				q			<=			16'h0381;
		end
		32'h0000D0C8: begin
				q			<=			16'h2C23;
		end
		32'h0000D0CA: begin
				q			<=			16'h04F1;
		end
		32'h0000D0CC: begin
				q			<=			16'h2783;
		end
		32'h0000D0CE: begin
				q			<=			16'h03C1;
		end
		32'h0000D0D0: begin
				q			<=			16'h2E23;
		end
		32'h0000D0D2: begin
				q			<=			16'h04F1;
		end
		32'h0000D0D4: begin
				q			<=			16'h0793;
		end
		32'h0000D0D6: begin
				q			<=			16'h0020;
		end
		32'h0000D0D8: begin
				q			<=			16'h8063;
		end
		32'h0000D0DA: begin
				q			<=			16'h28FB;
		end
		32'h0000D0DC: begin
				q			<=			16'h0793;
		end
		32'h0000D0DE: begin
				q			<=			16'h0030;
		end
		32'h0000D0E0: begin
				q			<=			16'h8A63;
		end
		32'h0000D0E2: begin
				q			<=			16'h28FB;
		end
		32'h0000D0E4: begin
				q			<=			16'h0793;
		end
		32'h0000D0E6: begin
				q			<=			16'h0010;
		end
		32'h0000D0E8: begin
				q			<=			16'h98E3;
		end
		32'h0000D0EA: begin
				q			<=			16'hE4FB;
		end
		32'h0000D0EC: begin
				q			<=			16'h2E23;
		end
		32'h0000D0EE: begin
				q			<=			16'h0401;
		end
		32'h0000D0F0: begin
				q			<=			16'h2C23;
		end
		32'h0000D0F2: begin
				q			<=			16'h0401;
		end
		32'h0000D0F4: begin
				q			<=			16'h2A23;
		end
		32'h0000D0F6: begin
				q			<=			16'h0401;
		end
		32'h0000D0F8: begin
				q			<=			16'h2823;
		end
		32'h0000D0FA: begin
				q			<=			16'h0401;
		end
		32'h0000D0FC: begin
				q			<=			16'h006F;
		end
		32'h0000D0FE: begin
				q			<=			16'h21C0;
		end
		32'h0000D100: begin
				q			<=			16'h2823;
		end
		32'h0000D102: begin
				q			<=			16'h0121;
		end
		32'h0000D104: begin
				q			<=			16'h2783;
		end
		32'h0000D106: begin
				q			<=			16'h0401;
		end
		32'h0000D108: begin
				q			<=			16'h0B93;
		end
		32'h0000D10A: begin
				q			<=			16'h0007;
		end
		32'h0000D10C: begin
				q			<=			16'h2823;
		end
		32'h0000D10E: begin
				q			<=			16'h04F1;
		end
		32'h0000D110: begin
				q			<=			16'h2783;
		end
		32'h0000D112: begin
				q			<=			16'h0441;
		end
		32'h0000D114: begin
				q			<=			16'h2A23;
		end
		32'h0000D116: begin
				q			<=			16'h04F1;
		end
		32'h0000D118: begin
				q			<=			16'h2783;
		end
		32'h0000D11A: begin
				q			<=			16'h0481;
		end
		32'h0000D11C: begin
				q			<=			16'h2C23;
		end
		32'h0000D11E: begin
				q			<=			16'h04F1;
		end
		32'h0000D120: begin
				q			<=			16'h2783;
		end
		32'h0000D122: begin
				q			<=			16'h04C1;
		end
		32'h0000D124: begin
				q			<=			16'h2E23;
		end
		32'h0000D126: begin
				q			<=			16'h04F1;
		end
		32'h0000D128: begin
				q			<=			16'hF06F;
		end
		32'h0000D12A: begin
				q			<=			16'hFADF;
		end
		32'h0000D12C: begin
				q			<=			16'h2783;
		end
		32'h0000D12E: begin
				q			<=			16'h0201;
		end
		32'h0000D130: begin
				q			<=			16'h2E23;
		end
		32'h0000D132: begin
				q			<=			16'h00F1;
		end
		32'h0000D134: begin
				q			<=			16'hF06F;
		end
		32'h0000D136: begin
				q			<=			16'hE05F;
		end
		32'h0000D138: begin
				q			<=			16'h2E23;
		end
		32'h0000D13A: begin
				q			<=			16'h0401;
		end
		32'h0000D13C: begin
				q			<=			16'h2C23;
		end
		32'h0000D13E: begin
				q			<=			16'h0401;
		end
		32'h0000D140: begin
				q			<=			16'h2A23;
		end
		32'h0000D142: begin
				q			<=			16'h0401;
		end
		32'h0000D144: begin
				q			<=			16'h2823;
		end
		32'h0000D146: begin
				q			<=			16'h0401;
		end
		32'h0000D148: begin
				q			<=			16'h0793;
		end
		32'h0000D14A: begin
				q			<=			16'hFFF7;
		end
		32'h0000D14C: begin
				q			<=			16'hF06F;
		end
		32'h0000D14E: begin
				q			<=			16'hEC1F;
		end
		32'h0000D150: begin
				q			<=			16'h0693;
		end
		32'h0000D152: begin
				q			<=			16'h0010;
		end
		32'h0000D154: begin
				q			<=			16'h87B3;
		end
		32'h0000D156: begin
				q			<=			16'h40F6;
		end
		32'h0000D158: begin
				q			<=			16'h0713;
		end
		32'h0000D15A: begin
				q			<=			16'h0740;
		end
		32'h0000D15C: begin
				q			<=			16'h4263;
		end
		32'h0000D15E: begin
				q			<=			16'h1CF7;
		end
		32'h0000D160: begin
				q			<=			16'hD613;
		end
		32'h0000D162: begin
				q			<=			16'h4057;
		end
		32'h0000D164: begin
				q			<=			16'hF693;
		end
		32'h0000D166: begin
				q			<=			16'h01F7;
		end
		32'h0000D168: begin
				q			<=			16'h0713;
		end
		32'h0000D16A: begin
				q			<=			16'h0000;
		end
		32'h0000D16C: begin
				q			<=			16'h0793;
		end
		32'h0000D16E: begin
				q			<=			16'h0000;
		end
		32'h0000D170: begin
				q			<=			16'h1593;
		end
		32'h0000D172: begin
				q			<=			16'h0027;
		end
		32'h0000D174: begin
				q			<=			16'h1263;
		end
		32'h0000D176: begin
				q			<=			16'h0AC7;
		end
		32'h0000D178: begin
				q			<=			16'h9863;
		end
		32'h0000D17A: begin
				q			<=			16'h0C06;
		end
		32'h0000D17C: begin
				q			<=			16'h0513;
		end
		32'h0000D17E: begin
				q			<=			16'h0030;
		end
		32'h0000D180: begin
				q			<=			16'h0613;
		end
		32'h0000D182: begin
				q			<=			16'h0501;
		end
		32'h0000D184: begin
				q			<=			16'h0533;
		end
		32'h0000D186: begin
				q			<=			16'h40E5;
		end
		32'h0000D188: begin
				q			<=			16'h5463;
		end
		32'h0000D18A: begin
				q			<=			16'h0AD5;
		end
		32'h0000D18C: begin
				q			<=			16'h0693;
		end
		32'h0000D18E: begin
				q			<=			16'h0040;
		end
		32'h0000D190: begin
				q			<=			16'h8733;
		end
		32'h0000D192: begin
				q			<=			16'h40E6;
		end
		32'h0000D194: begin
				q			<=			16'h0613;
		end
		32'h0000D196: begin
				q			<=			16'h0040;
		end
		32'h0000D198: begin
				q			<=			16'h1663;
		end
		32'h0000D19A: begin
				q			<=			16'h12C7;
		end
		32'h0000D19C: begin
				q			<=			16'h2683;
		end
		32'h0000D19E: begin
				q			<=			16'h0501;
		end
		32'h0000D1A0: begin
				q			<=			16'h37B3;
		end
		32'h0000D1A2: begin
				q			<=			16'h00F0;
		end
		32'h0000D1A4: begin
				q			<=			16'hE7B3;
		end
		32'h0000D1A6: begin
				q			<=			16'h00D7;
		end
		32'h0000D1A8: begin
				q			<=			16'h2823;
		end
		32'h0000D1AA: begin
				q			<=			16'h04F1;
		end
		32'h0000D1AC: begin
				q			<=			16'hF693;
		end
		32'h0000D1AE: begin
				q			<=			16'h0077;
		end
		32'h0000D1B0: begin
				q			<=			16'h8263;
		end
		32'h0000D1B2: begin
				q			<=			16'h0406;
		end
		32'h0000D1B4: begin
				q			<=			16'hF693;
		end
		32'h0000D1B6: begin
				q			<=			16'h00F7;
		end
		32'h0000D1B8: begin
				q			<=			16'h8E63;
		end
		32'h0000D1BA: begin
				q			<=			16'h02E6;
		end
		32'h0000D1BC: begin
				q			<=			16'h2703;
		end
		32'h0000D1BE: begin
				q			<=			16'h0541;
		end
		32'h0000D1C0: begin
				q			<=			16'h8793;
		end
		32'h0000D1C2: begin
				q			<=			16'h0047;
		end
		32'h0000D1C4: begin
				q			<=			16'h2823;
		end
		32'h0000D1C6: begin
				q			<=			16'h04F1;
		end
		32'h0000D1C8: begin
				q			<=			16'hB793;
		end
		32'h0000D1CA: begin
				q			<=			16'h0047;
		end
		32'h0000D1CC: begin
				q			<=			16'h8733;
		end
		32'h0000D1CE: begin
				q			<=			16'h00E7;
		end
		32'h0000D1D0: begin
				q			<=			16'h37B3;
		end
		32'h0000D1D2: begin
				q			<=			16'h00F7;
		end
		32'h0000D1D4: begin
				q			<=			16'h2A23;
		end
		32'h0000D1D6: begin
				q			<=			16'h04E1;
		end
		32'h0000D1D8: begin
				q			<=			16'h2703;
		end
		32'h0000D1DA: begin
				q			<=			16'h0581;
		end
		32'h0000D1DC: begin
				q			<=			16'h8733;
		end
		32'h0000D1DE: begin
				q			<=			16'h00E7;
		end
		32'h0000D1E0: begin
				q			<=			16'h2C23;
		end
		32'h0000D1E2: begin
				q			<=			16'h04E1;
		end
		32'h0000D1E4: begin
				q			<=			16'h3733;
		end
		32'h0000D1E6: begin
				q			<=			16'h00F7;
		end
		32'h0000D1E8: begin
				q			<=			16'h2783;
		end
		32'h0000D1EA: begin
				q			<=			16'h05C1;
		end
		32'h0000D1EC: begin
				q			<=			16'h0733;
		end
		32'h0000D1EE: begin
				q			<=			16'h00F7;
		end
		32'h0000D1F0: begin
				q			<=			16'h2E23;
		end
		32'h0000D1F2: begin
				q			<=			16'h04E1;
		end
		32'h0000D1F4: begin
				q			<=			16'h2783;
		end
		32'h0000D1F6: begin
				q			<=			16'h05C1;
		end
		32'h0000D1F8: begin
				q			<=			16'h9713;
		end
		32'h0000D1FA: begin
				q			<=			16'h00C7;
		end
		32'h0000D1FC: begin
				q			<=			16'h5063;
		end
		32'h0000D1FE: begin
				q			<=			16'h0E07;
		end
		32'h0000D200: begin
				q			<=			16'h2E23;
		end
		32'h0000D202: begin
				q			<=			16'h0401;
		end
		32'h0000D204: begin
				q			<=			16'h2C23;
		end
		32'h0000D206: begin
				q			<=			16'h0401;
		end
		32'h0000D208: begin
				q			<=			16'h2A23;
		end
		32'h0000D20A: begin
				q			<=			16'h0401;
		end
		32'h0000D20C: begin
				q			<=			16'h2823;
		end
		32'h0000D20E: begin
				q			<=			16'h0401;
		end
		32'h0000D210: begin
				q			<=			16'h0793;
		end
		32'h0000D212: begin
				q			<=			16'h0010;
		end
		32'h0000D214: begin
				q			<=			16'hF06F;
		end
		32'h0000D216: begin
				q			<=			16'hDF9F;
		end
		32'h0000D218: begin
				q			<=			16'h0513;
		end
		32'h0000D21A: begin
				q			<=			16'h0501;
		end
		32'h0000D21C: begin
				q			<=			16'h05B3;
		end
		32'h0000D21E: begin
				q			<=			16'h00B5;
		end
		32'h0000D220: begin
				q			<=			16'hA583;
		end
		32'h0000D222: begin
				q			<=			16'h0005;
		end
		32'h0000D224: begin
				q			<=			16'h0713;
		end
		32'h0000D226: begin
				q			<=			16'h0017;
		end
		32'h0000D228: begin
				q			<=			16'hE7B3;
		end
		32'h0000D22A: begin
				q			<=			16'h00B7;
		end
		32'h0000D22C: begin
				q			<=			16'hF06F;
		end
		32'h0000D22E: begin
				q			<=			16'hF45F;
		end
		32'h0000D230: begin
				q			<=			16'h0833;
		end
		32'h0000D232: begin
				q			<=			16'h00B6;
		end
		32'h0000D234: begin
				q			<=			16'h2803;
		end
		32'h0000D236: begin
				q			<=			16'h0008;
		end
		32'h0000D238: begin
				q			<=			16'h8693;
		end
		32'h0000D23A: begin
				q			<=			16'h0016;
		end
		32'h0000D23C: begin
				q			<=			16'h0613;
		end
		32'h0000D23E: begin
				q			<=			16'h0046;
		end
		32'h0000D240: begin
				q			<=			16'h2E23;
		end
		32'h0000D242: begin
				q			<=			16'hFF06;
		end
		32'h0000D244: begin
				q			<=			16'hF06F;
		end
		32'h0000D246: begin
				q			<=			16'hF45F;
		end
		32'h0000D248: begin
				q			<=			16'h0613;
		end
		32'h0000D24A: begin
				q			<=			16'h0801;
		end
		32'h0000D24C: begin
				q			<=			16'h0633;
		end
		32'h0000D24E: begin
				q			<=			16'h00B6;
		end
		32'h0000D250: begin
				q			<=			16'h2603;
		end
		32'h0000D252: begin
				q			<=			16'hFD06;
		end
		32'h0000D254: begin
				q			<=			16'h0813;
		end
		32'h0000D256: begin
				q			<=			16'h0200;
		end
		32'h0000D258: begin
				q			<=			16'h0833;
		end
		32'h0000D25A: begin
				q			<=			16'h40D8;
		end
		32'h0000D25C: begin
				q			<=			16'h1633;
		end
		32'h0000D25E: begin
				q			<=			16'h0106;
		end
		32'h0000D260: begin
				q			<=			16'hE7B3;
		end
		32'h0000D262: begin
				q			<=			16'h00C7;
		end
		32'h0000D264: begin
				q			<=			16'h0613;
		end
		32'h0000D266: begin
				q			<=			16'h0030;
		end
		32'h0000D268: begin
				q			<=			16'h0893;
		end
		32'h0000D26A: begin
				q			<=			16'h0501;
		end
		32'h0000D26C: begin
				q			<=			16'h0313;
		end
		32'h0000D26E: begin
				q			<=			16'h0000;
		end
		32'h0000D270: begin
				q			<=			16'h0633;
		end
		32'h0000D272: begin
				q			<=			16'h40E6;
		end
		32'h0000D274: begin
				q			<=			16'h4463;
		end
		32'h0000D276: begin
				q			<=			16'h02C3;
		end
		32'h0000D278: begin
				q			<=			16'h0593;
		end
		32'h0000D27A: begin
				q			<=			16'h0040;
		end
		32'h0000D27C: begin
				q			<=			16'h8733;
		end
		32'h0000D27E: begin
				q			<=			16'h40E5;
		end
		32'h0000D280: begin
				q			<=			16'h1613;
		end
		32'h0000D282: begin
				q			<=			16'h0026;
		end
		32'h0000D284: begin
				q			<=			16'h0593;
		end
		32'h0000D286: begin
				q			<=			16'h0801;
		end
		32'h0000D288: begin
				q			<=			16'h8633;
		end
		32'h0000D28A: begin
				q			<=			16'h00C5;
		end
		32'h0000D28C: begin
				q			<=			16'h2583;
		end
		32'h0000D28E: begin
				q			<=			16'h05C1;
		end
		32'h0000D290: begin
				q			<=			16'hD6B3;
		end
		32'h0000D292: begin
				q			<=			16'h00D5;
		end
		32'h0000D294: begin
				q			<=			16'h2823;
		end
		32'h0000D296: begin
				q			<=			16'hFCD6;
		end
		32'h0000D298: begin
				q			<=			16'hF06F;
		end
		32'h0000D29A: begin
				q			<=			16'hEFDF;
		end
		32'h0000D29C: begin
				q			<=			16'h8E33;
		end
		32'h0000D29E: begin
				q			<=			16'h00B8;
		end
		32'h0000D2A0: begin
				q			<=			16'h2503;
		end
		32'h0000D2A2: begin
				q			<=			16'h000E;
		end
		32'h0000D2A4: begin
				q			<=			16'h2E03;
		end
		32'h0000D2A6: begin
				q			<=			16'h004E;
		end
		32'h0000D2A8: begin
				q			<=			16'h0313;
		end
		32'h0000D2AA: begin
				q			<=			16'h0013;
		end
		32'h0000D2AC: begin
				q			<=			16'h5533;
		end
		32'h0000D2AE: begin
				q			<=			16'h00D5;
		end
		32'h0000D2B0: begin
				q			<=			16'h1E33;
		end
		32'h0000D2B2: begin
				q			<=			16'h010E;
		end
		32'h0000D2B4: begin
				q			<=			16'h6533;
		end
		32'h0000D2B6: begin
				q			<=			16'h01C5;
		end
		32'h0000D2B8: begin
				q			<=			16'hA023;
		end
		32'h0000D2BA: begin
				q			<=			16'h00A8;
		end
		32'h0000D2BC: begin
				q			<=			16'h8893;
		end
		32'h0000D2BE: begin
				q			<=			16'h0048;
		end
		32'h0000D2C0: begin
				q			<=			16'hF06F;
		end
		32'h0000D2C2: begin
				q			<=			16'hFB5F;
		end
		32'h0000D2C4: begin
				q			<=			16'h1693;
		end
		32'h0000D2C6: begin
				q			<=			16'h0027;
		end
		32'h0000D2C8: begin
				q			<=			16'h0593;
		end
		32'h0000D2CA: begin
				q			<=			16'h0501;
		end
		32'h0000D2CC: begin
				q			<=			16'h86B3;
		end
		32'h0000D2CE: begin
				q			<=			16'h00D5;
		end
		32'h0000D2D0: begin
				q			<=			16'hA023;
		end
		32'h0000D2D2: begin
				q			<=			16'h0006;
		end
		32'h0000D2D4: begin
				q			<=			16'h0713;
		end
		32'h0000D2D6: begin
				q			<=			16'h0017;
		end
		32'h0000D2D8: begin
				q			<=			16'hF06F;
		end
		32'h0000D2DA: begin
				q			<=			16'hEC1F;
		end
		32'h0000D2DC: begin
				q			<=			16'h0793;
		end
		32'h0000D2DE: begin
				q			<=			16'h0501;
		end
		32'h0000D2E0: begin
				q			<=			16'h0693;
		end
		32'h0000D2E2: begin
				q			<=			16'h0000;
		end
		32'h0000D2E4: begin
				q			<=			16'h0593;
		end
		32'h0000D2E6: begin
				q			<=			16'h0030;
		end
		32'h0000D2E8: begin
				q			<=			16'hA703;
		end
		32'h0000D2EA: begin
				q			<=			16'h0007;
		end
		32'h0000D2EC: begin
				q			<=			16'hA603;
		end
		32'h0000D2EE: begin
				q			<=			16'h0047;
		end
		32'h0000D2F0: begin
				q			<=			16'h8693;
		end
		32'h0000D2F2: begin
				q			<=			16'h0016;
		end
		32'h0000D2F4: begin
				q			<=			16'h5713;
		end
		32'h0000D2F6: begin
				q			<=			16'h0037;
		end
		32'h0000D2F8: begin
				q			<=			16'h1613;
		end
		32'h0000D2FA: begin
				q			<=			16'h01D6;
		end
		32'h0000D2FC: begin
				q			<=			16'h6733;
		end
		32'h0000D2FE: begin
				q			<=			16'h00C7;
		end
		32'h0000D300: begin
				q			<=			16'hA023;
		end
		32'h0000D302: begin
				q			<=			16'h00E7;
		end
		32'h0000D304: begin
				q			<=			16'h8793;
		end
		32'h0000D306: begin
				q			<=			16'h0047;
		end
		32'h0000D308: begin
				q			<=			16'h90E3;
		end
		32'h0000D30A: begin
				q			<=			16'hFEB6;
		end
		32'h0000D30C: begin
				q			<=			16'h2783;
		end
		32'h0000D30E: begin
				q			<=			16'h05C1;
		end
		32'h0000D310: begin
				q			<=			16'hD793;
		end
		32'h0000D312: begin
				q			<=			16'h0037;
		end
		32'h0000D314: begin
				q			<=			16'h2E23;
		end
		32'h0000D316: begin
				q			<=			16'h04F1;
		end
		32'h0000D318: begin
				q			<=			16'h0793;
		end
		32'h0000D31A: begin
				q			<=			16'h0000;
		end
		32'h0000D31C: begin
				q			<=			16'hF06F;
		end
		32'h0000D31E: begin
				q			<=			16'hCF1F;
		end
		32'h0000D320: begin
				q			<=			16'h2783;
		end
		32'h0000D322: begin
				q			<=			16'h0541;
		end
		32'h0000D324: begin
				q			<=			16'h2703;
		end
		32'h0000D326: begin
				q			<=			16'h0501;
		end
		32'h0000D328: begin
				q			<=			16'h6733;
		end
		32'h0000D32A: begin
				q			<=			16'h00F7;
		end
		32'h0000D32C: begin
				q			<=			16'h2783;
		end
		32'h0000D32E: begin
				q			<=			16'h0581;
		end
		32'h0000D330: begin
				q			<=			16'h6733;
		end
		32'h0000D332: begin
				q			<=			16'h00F7;
		end
		32'h0000D334: begin
				q			<=			16'h2783;
		end
		32'h0000D336: begin
				q			<=			16'h05C1;
		end
		32'h0000D338: begin
				q			<=			16'h6733;
		end
		32'h0000D33A: begin
				q			<=			16'h00F7;
		end
		32'h0000D33C: begin
				q			<=			16'h0793;
		end
		32'h0000D33E: begin
				q			<=			16'h0000;
		end
		32'h0000D340: begin
				q			<=			16'h06E3;
		end
		32'h0000D342: begin
				q			<=			16'hCC07;
		end
		32'h0000D344: begin
				q			<=			16'h2E23;
		end
		32'h0000D346: begin
				q			<=			16'h0401;
		end
		32'h0000D348: begin
				q			<=			16'h2C23;
		end
		32'h0000D34A: begin
				q			<=			16'h0401;
		end
		32'h0000D34C: begin
				q			<=			16'h2A23;
		end
		32'h0000D34E: begin
				q			<=			16'h0401;
		end
		32'h0000D350: begin
				q			<=			16'h2823;
		end
		32'h0000D352: begin
				q			<=			16'h0401;
		end
		32'h0000D354: begin
				q			<=			16'hF06F;
		end
		32'h0000D356: begin
				q			<=			16'hCB9F;
		end
		32'h0000D358: begin
				q			<=			16'h87B7;
		end
		32'h0000D35A: begin
				q			<=			16'h0000;
		end
		32'h0000D35C: begin
				q			<=			16'h2E23;
		end
		32'h0000D35E: begin
				q			<=			16'h0401;
		end
		32'h0000D360: begin
				q			<=			16'h2C23;
		end
		32'h0000D362: begin
				q			<=			16'h0401;
		end
		32'h0000D364: begin
				q			<=			16'h2A23;
		end
		32'h0000D366: begin
				q			<=			16'h0401;
		end
		32'h0000D368: begin
				q			<=			16'h2823;
		end
		32'h0000D36A: begin
				q			<=			16'h0401;
		end
		32'h0000D36C: begin
				q			<=			16'h8793;
		end
		32'h0000D36E: begin
				q			<=			16'hFFF7;
		end
		32'h0000D370: begin
				q			<=			16'hF06F;
		end
		32'h0000D372: begin
				q			<=			16'hC9DF;
		end
		32'h0000D374: begin
				q			<=			16'h87B7;
		end
		32'h0000D376: begin
				q			<=			16'h0000;
		end
		32'h0000D378: begin
				q			<=			16'h2E23;
		end
		32'h0000D37A: begin
				q			<=			16'h04F1;
		end
		32'h0000D37C: begin
				q			<=			16'h2C23;
		end
		32'h0000D37E: begin
				q			<=			16'h0401;
		end
		32'h0000D380: begin
				q			<=			16'h2A23;
		end
		32'h0000D382: begin
				q			<=			16'h0401;
		end
		32'h0000D384: begin
				q			<=			16'h2823;
		end
		32'h0000D386: begin
				q			<=			16'h0401;
		end
		32'h0000D388: begin
				q			<=			16'h8793;
		end
		32'h0000D38A: begin
				q			<=			16'hFFF7;
		end
		32'h0000D38C: begin
				q			<=			16'h2823;
		end
		32'h0000D38E: begin
				q			<=			16'h0001;
		end
		32'h0000D390: begin
				q			<=			16'hF06F;
		end
		32'h0000D392: begin
				q			<=			16'hC7DF;
		end
		32'h0000D394: begin
				q			<=			16'h0000;
		end
		32'h0000D396: begin
				q			<=			16'h0000;
		end
		32'h0000D398: begin
				q			<=			16'h0113;
		end
		32'h0000D39A: begin
				q			<=			16'hFA01;
		end
		32'h0000D39C: begin
				q			<=			16'hA783;
		end
		32'h0000D39E: begin
				q			<=			16'h0085;
		end
		32'h0000D3A0: begin
				q			<=			16'h2823;
		end
		32'h0000D3A2: begin
				q			<=			16'h0521;
		end
		32'h0000D3A4: begin
				q			<=			16'hA903;
		end
		32'h0000D3A6: begin
				q			<=			16'h00C5;
		end
		32'h0000D3A8: begin
				q			<=			16'hA683;
		end
		32'h0000D3AA: begin
				q			<=			16'h0005;
		end
		32'h0000D3AC: begin
				q			<=			16'hA703;
		end
		32'h0000D3AE: begin
				q			<=			16'h0045;
		end
		32'h0000D3B0: begin
				q			<=			16'h2A23;
		end
		32'h0000D3B2: begin
				q			<=			16'h0491;
		end
		32'h0000D3B4: begin
				q			<=			16'h2C23;
		end
		32'h0000D3B6: begin
				q			<=			16'h02F1;
		end
		32'h0000D3B8: begin
				q			<=			16'h0493;
		end
		32'h0000D3BA: begin
				q			<=			16'h0005;
		end
		32'h0000D3BC: begin
				q			<=			16'h2C23;
		end
		32'h0000D3BE: begin
				q			<=			16'h00F1;
		end
		32'h0000D3C0: begin
				q			<=			16'h2E03;
		end
		32'h0000D3C2: begin
				q			<=			16'h0006;
		end
		32'h0000D3C4: begin
				q			<=			16'h1793;
		end
		32'h0000D3C6: begin
				q			<=			16'h0109;
		end
		32'h0000D3C8: begin
				q			<=			16'h2303;
		end
		32'h0000D3CA: begin
				q			<=			16'h0046;
		end
		32'h0000D3CC: begin
				q			<=			16'h2883;
		end
		32'h0000D3CE: begin
				q			<=			16'h0086;
		end
		32'h0000D3D0: begin
				q			<=			16'h2503;
		end
		32'h0000D3D2: begin
				q			<=			16'h00C6;
		end
		32'h0000D3D4: begin
				q			<=			16'h2C23;
		end
		32'h0000D3D6: begin
				q			<=			16'h0481;
		end
		32'h0000D3D8: begin
				q			<=			16'hD793;
		end
		32'h0000D3DA: begin
				q			<=			16'h0107;
		end
		32'h0000D3DC: begin
				q			<=			16'h1413;
		end
		32'h0000D3DE: begin
				q			<=			16'h0019;
		end
		32'h0000D3E0: begin
				q			<=			16'h2E23;
		end
		32'h0000D3E2: begin
				q			<=			16'h0321;
		end
		32'h0000D3E4: begin
				q			<=			16'h2E23;
		end
		32'h0000D3E6: begin
				q			<=			16'h0411;
		end
		32'h0000D3E8: begin
				q			<=			16'h2623;
		end
		32'h0000D3EA: begin
				q			<=			16'h0531;
		end
		32'h0000D3EC: begin
				q			<=			16'h2423;
		end
		32'h0000D3EE: begin
				q			<=			16'h0541;
		end
		32'h0000D3F0: begin
				q			<=			16'h2223;
		end
		32'h0000D3F2: begin
				q			<=			16'h0551;
		end
		32'h0000D3F4: begin
				q			<=			16'h2823;
		end
		32'h0000D3F6: begin
				q			<=			16'h02D1;
		end
		32'h0000D3F8: begin
				q			<=			16'h2A23;
		end
		32'h0000D3FA: begin
				q			<=			16'h02E1;
		end
		32'h0000D3FC: begin
				q			<=			16'h2823;
		end
		32'h0000D3FE: begin
				q			<=			16'h00D1;
		end
		32'h0000D400: begin
				q			<=			16'h2A23;
		end
		32'h0000D402: begin
				q			<=			16'h00E1;
		end
		32'h0000D404: begin
				q			<=			16'h2E23;
		end
		32'h0000D406: begin
				q			<=			16'h00F1;
		end
		32'h0000D408: begin
				q			<=			16'h5413;
		end
		32'h0000D40A: begin
				q			<=			16'h0114;
		end
		32'h0000D40C: begin
				q			<=			16'h5913;
		end
		32'h0000D40E: begin
				q			<=			16'h01F9;
		end
		32'h0000D410: begin
				q			<=			16'h0813;
		end
		32'h0000D412: begin
				q			<=			16'h0101;
		end
		32'h0000D414: begin
				q			<=			16'h0593;
		end
		32'h0000D416: begin
				q			<=			16'h01C1;
		end
		32'h0000D418: begin
				q			<=			16'hA783;
		end
		32'h0000D41A: begin
				q			<=			16'h0005;
		end
		32'h0000D41C: begin
				q			<=			16'hA703;
		end
		32'h0000D41E: begin
				q			<=			16'hFFC5;
		end
		32'h0000D420: begin
				q			<=			16'h8593;
		end
		32'h0000D422: begin
				q			<=			16'hFFC5;
		end
		32'h0000D424: begin
				q			<=			16'h9793;
		end
		32'h0000D426: begin
				q			<=			16'h0037;
		end
		32'h0000D428: begin
				q			<=			16'h5713;
		end
		32'h0000D42A: begin
				q			<=			16'h01D7;
		end
		32'h0000D42C: begin
				q			<=			16'hE7B3;
		end
		32'h0000D42E: begin
				q			<=			16'h00E7;
		end
		32'h0000D430: begin
				q			<=			16'hA223;
		end
		32'h0000D432: begin
				q			<=			16'h00F5;
		end
		32'h0000D434: begin
				q			<=			16'h12E3;
		end
		32'h0000D436: begin
				q			<=			16'hFEB8;
		end
		32'h0000D438: begin
				q			<=			16'h2683;
		end
		32'h0000D43A: begin
				q			<=			16'h0101;
		end
		32'h0000D43C: begin
				q			<=			16'h1793;
		end
		32'h0000D43E: begin
				q			<=			16'h0105;
		end
		32'h0000D440: begin
				q			<=			16'h1613;
		end
		32'h0000D442: begin
				q			<=			16'h0015;
		end
		32'h0000D444: begin
				q			<=			16'h9693;
		end
		32'h0000D446: begin
				q			<=			16'h0036;
		end
		32'h0000D448: begin
				q			<=			16'hD793;
		end
		32'h0000D44A: begin
				q			<=			16'h0107;
		end
		32'h0000D44C: begin
				q			<=			16'h2A23;
		end
		32'h0000D44E: begin
				q			<=			16'h0261;
		end
		32'h0000D450: begin
				q			<=			16'h2C23;
		end
		32'h0000D452: begin
				q			<=			16'h0311;
		end
		32'h0000D454: begin
				q			<=			16'h2E23;
		end
		32'h0000D456: begin
				q			<=			16'h02A1;
		end
		32'h0000D458: begin
				q			<=			16'h2223;
		end
		32'h0000D45A: begin
				q			<=			16'h0261;
		end
		32'h0000D45C: begin
				q			<=			16'h2423;
		end
		32'h0000D45E: begin
				q			<=			16'h0311;
		end
		32'h0000D460: begin
				q			<=			16'h2823;
		end
		32'h0000D462: begin
				q			<=			16'h00D1;
		end
		32'h0000D464: begin
				q			<=			16'h2823;
		end
		32'h0000D466: begin
				q			<=			16'h03C1;
		end
		32'h0000D468: begin
				q			<=			16'h2023;
		end
		32'h0000D46A: begin
				q			<=			16'h03C1;
		end
		32'h0000D46C: begin
				q			<=			16'h2623;
		end
		32'h0000D46E: begin
				q			<=			16'h02F1;
		end
		32'h0000D470: begin
				q			<=			16'h5613;
		end
		32'h0000D472: begin
				q			<=			16'h0116;
		end
		32'h0000D474: begin
				q			<=			16'h5513;
		end
		32'h0000D476: begin
				q			<=			16'h01F5;
		end
		32'h0000D478: begin
				q			<=			16'h0893;
		end
		32'h0000D47A: begin
				q			<=			16'h0201;
		end
		32'h0000D47C: begin
				q			<=			16'h0313;
		end
		32'h0000D47E: begin
				q			<=			16'h02C1;
		end
		32'h0000D480: begin
				q			<=			16'h2783;
		end
		32'h0000D482: begin
				q			<=			16'h0003;
		end
		32'h0000D484: begin
				q			<=			16'h2703;
		end
		32'h0000D486: begin
				q			<=			16'hFFC3;
		end
		32'h0000D488: begin
				q			<=			16'h0313;
		end
		32'h0000D48A: begin
				q			<=			16'hFFC3;
		end
		32'h0000D48C: begin
				q			<=			16'h9793;
		end
		32'h0000D48E: begin
				q			<=			16'h0037;
		end
		32'h0000D490: begin
				q			<=			16'h5713;
		end
		32'h0000D492: begin
				q			<=			16'h01D7;
		end
		32'h0000D494: begin
				q			<=			16'hE7B3;
		end
		32'h0000D496: begin
				q			<=			16'h00E7;
		end
		32'h0000D498: begin
				q			<=			16'h2223;
		end
		32'h0000D49A: begin
				q			<=			16'h00F3;
		end
		32'h0000D49C: begin
				q			<=			16'h92E3;
		end
		32'h0000D49E: begin
				q			<=			16'hFE68;
		end
		32'h0000D4A0: begin
				q			<=			16'h2783;
		end
		32'h0000D4A2: begin
				q			<=			16'h0201;
		end
		32'h0000D4A4: begin
				q			<=			16'h8737;
		end
		32'h0000D4A6: begin
				q			<=			16'h0000;
		end
		32'h0000D4A8: begin
				q			<=			16'h0713;
		end
		32'h0000D4AA: begin
				q			<=			16'hFFF7;
		end
		32'h0000D4AC: begin
				q			<=			16'h9793;
		end
		32'h0000D4AE: begin
				q			<=			16'h0037;
		end
		32'h0000D4B0: begin
				q			<=			16'h2023;
		end
		32'h0000D4B2: begin
				q			<=			16'h02F1;
		end
		32'h0000D4B4: begin
				q			<=			16'h1063;
		end
		32'h0000D4B6: begin
				q			<=			16'h02E6;
		end
		32'h0000D4B8: begin
				q			<=			16'h2E03;
		end
		32'h0000D4BA: begin
				q			<=			16'h0281;
		end
		32'h0000D4BC: begin
				q			<=			16'h2703;
		end
		32'h0000D4BE: begin
				q			<=			16'h0241;
		end
		32'h0000D4C0: begin
				q			<=			16'h6733;
		end
		32'h0000D4C2: begin
				q			<=			16'h01C7;
		end
		32'h0000D4C4: begin
				q			<=			16'h2E03;
		end
		32'h0000D4C6: begin
				q			<=			16'h02C1;
		end
		32'h0000D4C8: begin
				q			<=			16'h6733;
		end
		32'h0000D4CA: begin
				q			<=			16'h01C7;
		end
		32'h0000D4CC: begin
				q			<=			16'h6733;
		end
		32'h0000D4CE: begin
				q			<=			16'h00F7;
		end
		32'h0000D4D0: begin
				q			<=			16'h1463;
		end
		32'h0000D4D2: begin
				q			<=			16'h0007;
		end
		32'h0000D4D4: begin
				q			<=			16'h4513;
		end
		32'h0000D4D6: begin
				q			<=			16'h0015;
		end
		32'h0000D4D8: begin
				q			<=			16'h0733;
		end
		32'h0000D4DA: begin
				q			<=			16'h40C4;
		end
		32'h0000D4DC: begin
				q			<=			16'h18E3;
		end
		32'h0000D4DE: begin
				q			<=			16'h1125;
		end
		32'h0000D4E0: begin
				q			<=			16'h5463;
		end
		32'h0000D4E2: begin
				q			<=			16'h30E0;
		end
		32'h0000D4E4: begin
				q			<=			16'h1863;
		end
		32'h0000D4E6: begin
				q			<=			16'h1406;
		end
		32'h0000D4E8: begin
				q			<=			16'h2503;
		end
		32'h0000D4EA: begin
				q			<=			16'h0241;
		end
		32'h0000D4EC: begin
				q			<=			16'h2583;
		end
		32'h0000D4EE: begin
				q			<=			16'h0281;
		end
		32'h0000D4F0: begin
				q			<=			16'h2803;
		end
		32'h0000D4F2: begin
				q			<=			16'h02C1;
		end
		32'h0000D4F4: begin
				q			<=			16'h6633;
		end
		32'h0000D4F6: begin
				q			<=			16'h00B5;
		end
		32'h0000D4F8: begin
				q			<=			16'h6633;
		end
		32'h0000D4FA: begin
				q			<=			16'h0106;
		end
		32'h0000D4FC: begin
				q			<=			16'h6633;
		end
		32'h0000D4FE: begin
				q			<=			16'h00F6;
		end
		32'h0000D500: begin
				q			<=			16'h1463;
		end
		32'h0000D502: begin
				q			<=			16'h0206;
		end
		32'h0000D504: begin
				q			<=			16'h2783;
		end
		32'h0000D506: begin
				q			<=			16'h0141;
		end
		32'h0000D508: begin
				q			<=			16'h2823;
		end
		32'h0000D50A: begin
				q			<=			16'h02D1;
		end
		32'h0000D50C: begin
				q			<=			16'h0413;
		end
		32'h0000D50E: begin
				q			<=			16'h0007;
		end
		32'h0000D510: begin
				q			<=			16'h2A23;
		end
		32'h0000D512: begin
				q			<=			16'h02F1;
		end
		32'h0000D514: begin
				q			<=			16'h2783;
		end
		32'h0000D516: begin
				q			<=			16'h0181;
		end
		32'h0000D518: begin
				q			<=			16'h2C23;
		end
		32'h0000D51A: begin
				q			<=			16'h02F1;
		end
		32'h0000D51C: begin
				q			<=			16'h2783;
		end
		32'h0000D51E: begin
				q			<=			16'h01C1;
		end
		32'h0000D520: begin
				q			<=			16'h2E23;
		end
		32'h0000D522: begin
				q			<=			16'h02F1;
		end
		32'h0000D524: begin
				q			<=			16'h006F;
		end
		32'h0000D526: begin
				q			<=			16'h3080;
		end
		32'h0000D528: begin
				q			<=			16'h0613;
		end
		32'h0000D52A: begin
				q			<=			16'hFFF7;
		end
		32'h0000D52C: begin
				q			<=			16'h1E63;
		end
		32'h0000D52E: begin
				q			<=			16'h0C06;
		end
		32'h0000D530: begin
				q			<=			16'h2703;
		end
		32'h0000D532: begin
				q			<=			16'h0141;
		end
		32'h0000D534: begin
				q			<=			16'h87B3;
		end
		32'h0000D536: begin
				q			<=			16'h00F6;
		end
		32'h0000D538: begin
				q			<=			16'hB6B3;
		end
		32'h0000D53A: begin
				q			<=			16'h00D7;
		end
		32'h0000D53C: begin
				q			<=			16'h0633;
		end
		32'h0000D53E: begin
				q			<=			16'h00E5;
		end
		32'h0000D540: begin
				q			<=			16'h2823;
		end
		32'h0000D542: begin
				q			<=			16'h02F1;
		end
		32'h0000D544: begin
				q			<=			16'h07B3;
		end
		32'h0000D546: begin
				q			<=			16'h00D6;
		end
		32'h0000D548: begin
				q			<=			16'hB6B3;
		end
		32'h0000D54A: begin
				q			<=			16'h00D7;
		end
		32'h0000D54C: begin
				q			<=			16'h2A23;
		end
		32'h0000D54E: begin
				q			<=			16'h02F1;
		end
		32'h0000D550: begin
				q			<=			16'h2783;
		end
		32'h0000D552: begin
				q			<=			16'h0181;
		end
		32'h0000D554: begin
				q			<=			16'h3733;
		end
		32'h0000D556: begin
				q			<=			16'h00E6;
		end
		32'h0000D558: begin
				q			<=			16'h66B3;
		end
		32'h0000D55A: begin
				q			<=			16'h00D7;
		end
		32'h0000D55C: begin
				q			<=			16'h8733;
		end
		32'h0000D55E: begin
				q			<=			16'h00F5;
		end
		32'h0000D560: begin
				q			<=			16'h0633;
		end
		32'h0000D562: begin
				q			<=			16'h00D7;
		end
		32'h0000D564: begin
				q			<=			16'h37B3;
		end
		32'h0000D566: begin
				q			<=			16'h00F7;
		end
		32'h0000D568: begin
				q			<=			16'h2703;
		end
		32'h0000D56A: begin
				q			<=			16'h01C1;
		end
		32'h0000D56C: begin
				q			<=			16'h36B3;
		end
		32'h0000D56E: begin
				q			<=			16'h00D6;
		end
		32'h0000D570: begin
				q			<=			16'hE7B3;
		end
		32'h0000D572: begin
				q			<=			16'h00D7;
		end
		32'h0000D574: begin
				q			<=			16'h0833;
		end
		32'h0000D576: begin
				q			<=			16'h00E8;
		end
		32'h0000D578: begin
				q			<=			16'h87B3;
		end
		32'h0000D57A: begin
				q			<=			16'h0107;
		end
		32'h0000D57C: begin
				q			<=			16'h2C23;
		end
		32'h0000D57E: begin
				q			<=			16'h02C1;
		end
		32'h0000D580: begin
				q			<=			16'h2E23;
		end
		32'h0000D582: begin
				q			<=			16'h02F1;
		end
		32'h0000D584: begin
				q			<=			16'h0413;
		end
		32'h0000D586: begin
				q			<=			16'h0010;
		end
		32'h0000D588: begin
				q			<=			16'h2783;
		end
		32'h0000D58A: begin
				q			<=			16'h03C1;
		end
		32'h0000D58C: begin
				q			<=			16'h9713;
		end
		32'h0000D58E: begin
				q			<=			16'h00C7;
		end
		32'h0000D590: begin
				q			<=			16'h5E63;
		end
		32'h0000D592: begin
				q			<=			16'h2807;
		end
		32'h0000D594: begin
				q			<=			16'h0737;
		end
		32'h0000D596: begin
				q			<=			16'hFFF8;
		end
		32'h0000D598: begin
				q			<=			16'h0713;
		end
		32'h0000D59A: begin
				q			<=			16'hFFF7;
		end
		32'h0000D59C: begin
				q			<=			16'hF7B3;
		end
		32'h0000D59E: begin
				q			<=			16'h00E7;
		end
		32'h0000D5A0: begin
				q			<=			16'h2E23;
		end
		32'h0000D5A2: begin
				q			<=			16'h02F1;
		end
		32'h0000D5A4: begin
				q			<=			16'h2783;
		end
		32'h0000D5A6: begin
				q			<=			16'h0301;
		end
		32'h0000D5A8: begin
				q			<=			16'h0413;
		end
		32'h0000D5AA: begin
				q			<=			16'h0014;
		end
		32'h0000D5AC: begin
				q			<=			16'h0713;
		end
		32'h0000D5AE: begin
				q			<=			16'h0301;
		end
		32'h0000D5B0: begin
				q			<=			16'h9793;
		end
		32'h0000D5B2: begin
				q			<=			16'h01F7;
		end
		32'h0000D5B4: begin
				q			<=			16'h0613;
		end
		32'h0000D5B6: begin
				q			<=			16'h0000;
		end
		32'h0000D5B8: begin
				q			<=			16'h0513;
		end
		32'h0000D5BA: begin
				q			<=			16'h0030;
		end
		32'h0000D5BC: begin
				q			<=			16'h2683;
		end
		32'h0000D5BE: begin
				q			<=			16'h0007;
		end
		32'h0000D5C0: begin
				q			<=			16'h2583;
		end
		32'h0000D5C2: begin
				q			<=			16'h0047;
		end
		32'h0000D5C4: begin
				q			<=			16'h0613;
		end
		32'h0000D5C6: begin
				q			<=			16'h0016;
		end
		32'h0000D5C8: begin
				q			<=			16'hD693;
		end
		32'h0000D5CA: begin
				q			<=			16'h0016;
		end
		32'h0000D5CC: begin
				q			<=			16'h9593;
		end
		32'h0000D5CE: begin
				q			<=			16'h01F5;
		end
		32'h0000D5D0: begin
				q			<=			16'hE6B3;
		end
		32'h0000D5D2: begin
				q			<=			16'h00B6;
		end
		32'h0000D5D4: begin
				q			<=			16'h2023;
		end
		32'h0000D5D6: begin
				q			<=			16'h00D7;
		end
		32'h0000D5D8: begin
				q			<=			16'h0713;
		end
		32'h0000D5DA: begin
				q			<=			16'h0047;
		end
		32'h0000D5DC: begin
				q			<=			16'h10E3;
		end
		32'h0000D5DE: begin
				q			<=			16'hFEA6;
		end
		32'h0000D5E0: begin
				q			<=			16'h2703;
		end
		32'h0000D5E2: begin
				q			<=			16'h03C1;
		end
		32'h0000D5E4: begin
				q			<=			16'h37B3;
		end
		32'h0000D5E6: begin
				q			<=			16'h00F0;
		end
		32'h0000D5E8: begin
				q			<=			16'h5713;
		end
		32'h0000D5EA: begin
				q			<=			16'h0017;
		end
		32'h0000D5EC: begin
				q			<=			16'h2E23;
		end
		32'h0000D5EE: begin
				q			<=			16'h02E1;
		end
		32'h0000D5F0: begin
				q			<=			16'h2703;
		end
		32'h0000D5F2: begin
				q			<=			16'h0301;
		end
		32'h0000D5F4: begin
				q			<=			16'h67B3;
		end
		32'h0000D5F6: begin
				q			<=			16'h00F7;
		end
		32'h0000D5F8: begin
				q			<=			16'h2823;
		end
		32'h0000D5FA: begin
				q			<=			16'h02F1;
		end
		32'h0000D5FC: begin
				q			<=			16'h87B7;
		end
		32'h0000D5FE: begin
				q			<=			16'h0000;
		end
		32'h0000D600: begin
				q			<=			16'h8793;
		end
		32'h0000D602: begin
				q			<=			16'hFFF7;
		end
		32'h0000D604: begin
				q			<=			16'h006F;
		end
		32'h0000D606: begin
				q			<=			16'h7D00;
		end
		32'h0000D608: begin
				q			<=			16'h87B7;
		end
		32'h0000D60A: begin
				q			<=			16'h0000;
		end
		32'h0000D60C: begin
				q			<=			16'h8793;
		end
		32'h0000D60E: begin
				q			<=			16'hFFF7;
		end
		32'h0000D610: begin
				q			<=			16'h0AE3;
		end
		32'h0000D612: begin
				q			<=			16'hEEF7;
		end
		32'h0000D614: begin
				q			<=			16'h0793;
		end
		32'h0000D616: begin
				q			<=			16'h0740;
		end
		32'h0000D618: begin
				q			<=			16'hD263;
		end
		32'h0000D61A: begin
				q			<=			16'h06C7;
		end
		32'h0000D61C: begin
				q			<=			16'h0793;
		end
		32'h0000D61E: begin
				q			<=			16'h0010;
		end
		32'h0000D620: begin
				q			<=			16'h2623;
		end
		32'h0000D622: begin
				q			<=			16'h0201;
		end
		32'h0000D624: begin
				q			<=			16'h2423;
		end
		32'h0000D626: begin
				q			<=			16'h0201;
		end
		32'h0000D628: begin
				q			<=			16'h2223;
		end
		32'h0000D62A: begin
				q			<=			16'h0201;
		end
		32'h0000D62C: begin
				q			<=			16'h2023;
		end
		32'h0000D62E: begin
				q			<=			16'h02F1;
		end
		32'h0000D630: begin
				q			<=			16'h006F;
		end
		32'h0000D632: begin
				q			<=			16'h0940;
		end
		32'h0000D634: begin
				q			<=			16'h87B7;
		end
		32'h0000D636: begin
				q			<=			16'h0000;
		end
		32'h0000D638: begin
				q			<=			16'h8793;
		end
		32'h0000D63A: begin
				q			<=			16'hFFF7;
		end
		32'h0000D63C: begin
				q			<=			16'h1263;
		end
		32'h0000D63E: begin
				q			<=			16'h02F4;
		end
		32'h0000D640: begin
				q			<=			16'h2783;
		end
		32'h0000D642: begin
				q			<=			16'h0141;
		end
		32'h0000D644: begin
				q			<=			16'h2823;
		end
		32'h0000D646: begin
				q			<=			16'h02D1;
		end
		32'h0000D648: begin
				q			<=			16'h2A23;
		end
		32'h0000D64A: begin
				q			<=			16'h02F1;
		end
		32'h0000D64C: begin
				q			<=			16'h2783;
		end
		32'h0000D64E: begin
				q			<=			16'h0181;
		end
		32'h0000D650: begin
				q			<=			16'h2C23;
		end
		32'h0000D652: begin
				q			<=			16'h02F1;
		end
		32'h0000D654: begin
				q			<=			16'h2783;
		end
		32'h0000D656: begin
				q			<=			16'h01C1;
		end
		32'h0000D658: begin
				q			<=			16'h2E23;
		end
		32'h0000D65A: begin
				q			<=			16'h02F1;
		end
		32'h0000D65C: begin
				q			<=			16'h006F;
		end
		32'h0000D65E: begin
				q			<=			16'h1D00;
		end
		32'h0000D660: begin
				q			<=			16'h2783;
		end
		32'h0000D662: begin
				q			<=			16'h02C1;
		end
		32'h0000D664: begin
				q			<=			16'h06B7;
		end
		32'h0000D666: begin
				q			<=			16'h0008;
		end
		32'h0000D668: begin
				q			<=			16'hE7B3;
		end
		32'h0000D66A: begin
				q			<=			16'h00D7;
		end
		32'h0000D66C: begin
				q			<=			16'h2623;
		end
		32'h0000D66E: begin
				q			<=			16'h02F1;
		end
		32'h0000D670: begin
				q			<=			16'h0793;
		end
		32'h0000D672: begin
				q			<=			16'h0740;
		end
		32'h0000D674: begin
				q			<=			16'hC4E3;
		end
		32'h0000D676: begin
				q			<=			16'hFAE7;
		end
		32'h0000D678: begin
				q			<=			16'h0613;
		end
		32'h0000D67A: begin
				q			<=			16'h0007;
		end
		32'h0000D67C: begin
				q			<=			16'h5693;
		end
		32'h0000D67E: begin
				q			<=			16'h4056;
		end
		32'h0000D680: begin
				q			<=			16'h7713;
		end
		32'h0000D682: begin
				q			<=			16'h01F6;
		end
		32'h0000D684: begin
				q			<=			16'h0793;
		end
		32'h0000D686: begin
				q			<=			16'h0000;
		end
		32'h0000D688: begin
				q			<=			16'h0613;
		end
		32'h0000D68A: begin
				q			<=			16'h0000;
		end
		32'h0000D68C: begin
				q			<=			16'h9593;
		end
		32'h0000D68E: begin
				q			<=			16'h0027;
		end
		32'h0000D690: begin
				q			<=			16'h9063;
		end
		32'h0000D692: begin
				q			<=			16'h0AD7;
		end
		32'h0000D694: begin
				q			<=			16'h1463;
		end
		32'h0000D696: begin
				q			<=			16'h0C07;
		end
		32'h0000D698: begin
				q			<=			16'h0693;
		end
		32'h0000D69A: begin
				q			<=			16'h0030;
		end
		32'h0000D69C: begin
				q			<=			16'h86B3;
		end
		32'h0000D69E: begin
				q			<=			16'h40F6;
		end
		32'h0000D6A0: begin
				q			<=			16'hD263;
		end
		32'h0000D6A2: begin
				q			<=			16'h0AE6;
		end
		32'h0000D6A4: begin
				q			<=			16'h0713;
		end
		32'h0000D6A6: begin
				q			<=			16'h0040;
		end
		32'h0000D6A8: begin
				q			<=			16'h07B3;
		end
		32'h0000D6AA: begin
				q			<=			16'h40F7;
		end
		32'h0000D6AC: begin
				q			<=			16'h0693;
		end
		32'h0000D6AE: begin
				q			<=			16'h0040;
		end
		32'h0000D6B0: begin
				q			<=			16'h9263;
		end
		32'h0000D6B2: begin
				q			<=			16'h12D7;
		end
		32'h0000D6B4: begin
				q			<=			16'h2783;
		end
		32'h0000D6B6: begin
				q			<=			16'h0201;
		end
		32'h0000D6B8: begin
				q			<=			16'h3633;
		end
		32'h0000D6BA: begin
				q			<=			16'h00C0;
		end
		32'h0000D6BC: begin
				q			<=			16'hE633;
		end
		32'h0000D6BE: begin
				q			<=			16'h00C7;
		end
		32'h0000D6C0: begin
				q			<=			16'h2023;
		end
		32'h0000D6C2: begin
				q			<=			16'h02C1;
		end
		32'h0000D6C4: begin
				q			<=			16'h2683;
		end
		32'h0000D6C6: begin
				q			<=			16'h0101;
		end
		32'h0000D6C8: begin
				q			<=			16'h2783;
		end
		32'h0000D6CA: begin
				q			<=			16'h0201;
		end
		32'h0000D6CC: begin
				q			<=			16'h2703;
		end
		32'h0000D6CE: begin
				q			<=			16'h0141;
		end
		32'h0000D6D0: begin
				q			<=			16'h2583;
		end
		32'h0000D6D2: begin
				q			<=			16'h0281;
		end
		32'h0000D6D4: begin
				q			<=			16'h87B3;
		end
		32'h0000D6D6: begin
				q			<=			16'h00F6;
		end
		32'h0000D6D8: begin
				q			<=			16'hB6B3;
		end
		32'h0000D6DA: begin
				q			<=			16'h00D7;
		end
		32'h0000D6DC: begin
				q			<=			16'h2823;
		end
		32'h0000D6DE: begin
				q			<=			16'h02F1;
		end
		32'h0000D6E0: begin
				q			<=			16'h2783;
		end
		32'h0000D6E2: begin
				q			<=			16'h0241;
		end
		32'h0000D6E4: begin
				q			<=			16'h2503;
		end
		32'h0000D6E6: begin
				q			<=			16'h02C1;
		end
		32'h0000D6E8: begin
				q			<=			16'h07B3;
		end
		32'h0000D6EA: begin
				q			<=			16'h00F7;
		end
		32'h0000D6EC: begin
				q			<=			16'h8633;
		end
		32'h0000D6EE: begin
				q			<=			16'h00D7;
		end
		32'h0000D6F0: begin
				q			<=			16'hB733;
		end
		32'h0000D6F2: begin
				q			<=			16'h00E7;
		end
		32'h0000D6F4: begin
				q			<=			16'h37B3;
		end
		32'h0000D6F6: begin
				q			<=			16'h00D6;
		end
		32'h0000D6F8: begin
				q			<=			16'h67B3;
		end
		32'h0000D6FA: begin
				q			<=			16'h00F7;
		end
		32'h0000D6FC: begin
				q			<=			16'h2703;
		end
		32'h0000D6FE: begin
				q			<=			16'h0181;
		end
		32'h0000D700: begin
				q			<=			16'h2683;
		end
		32'h0000D702: begin
				q			<=			16'h01C1;
		end
		32'h0000D704: begin
				q			<=			16'h2A23;
		end
		32'h0000D706: begin
				q			<=			16'h02C1;
		end
		32'h0000D708: begin
				q			<=			16'h05B3;
		end
		32'h0000D70A: begin
				q			<=			16'h00B7;
		end
		32'h0000D70C: begin
				q			<=			16'h8633;
		end
		32'h0000D70E: begin
				q			<=			16'h00F5;
		end
		32'h0000D710: begin
				q			<=			16'hB733;
		end
		32'h0000D712: begin
				q			<=			16'h00E5;
		end
		32'h0000D714: begin
				q			<=			16'h37B3;
		end
		32'h0000D716: begin
				q			<=			16'h00F6;
		end
		32'h0000D718: begin
				q			<=			16'h86B3;
		end
		32'h0000D71A: begin
				q			<=			16'h00A6;
		end
		32'h0000D71C: begin
				q			<=			16'h6733;
		end
		32'h0000D71E: begin
				q			<=			16'h00F7;
		end
		32'h0000D720: begin
				q			<=			16'h8733;
		end
		32'h0000D722: begin
				q			<=			16'h00E6;
		end
		32'h0000D724: begin
				q			<=			16'h2C23;
		end
		32'h0000D726: begin
				q			<=			16'h02C1;
		end
		32'h0000D728: begin
				q			<=			16'h2E23;
		end
		32'h0000D72A: begin
				q			<=			16'h02E1;
		end
		32'h0000D72C: begin
				q			<=			16'hF06F;
		end
		32'h0000D72E: begin
				q			<=			16'hE5DF;
		end
		32'h0000D730: begin
				q			<=			16'h85B3;
		end
		32'h0000D732: begin
				q			<=			16'h00B8;
		end
		32'h0000D734: begin
				q			<=			16'hA583;
		end
		32'h0000D736: begin
				q			<=			16'h0005;
		end
		32'h0000D738: begin
				q			<=			16'h8793;
		end
		32'h0000D73A: begin
				q			<=			16'h0017;
		end
		32'h0000D73C: begin
				q			<=			16'h6633;
		end
		32'h0000D73E: begin
				q			<=			16'h00B6;
		end
		32'h0000D740: begin
				q			<=			16'hF06F;
		end
		32'h0000D742: begin
				q			<=			16'hF4DF;
		end
		32'h0000D744: begin
				q			<=			16'h0533;
		end
		32'h0000D746: begin
				q			<=			16'h00B3;
		end
		32'h0000D748: begin
				q			<=			16'h2503;
		end
		32'h0000D74A: begin
				q			<=			16'h0005;
		end
		32'h0000D74C: begin
				q			<=			16'h0713;
		end
		32'h0000D74E: begin
				q			<=			16'h0017;
		end
		32'h0000D750: begin
				q			<=			16'h0313;
		end
		32'h0000D752: begin
				q			<=			16'h0043;
		end
		32'h0000D754: begin
				q			<=			16'h2E23;
		end
		32'h0000D756: begin
				q			<=			16'hFEA3;
		end
		32'h0000D758: begin
				q			<=			16'hF06F;
		end
		32'h0000D75A: begin
				q			<=			16'hF49F;
		end
		32'h0000D75C: begin
				q			<=			16'h0693;
		end
		32'h0000D75E: begin
				q			<=			16'h0401;
		end
		32'h0000D760: begin
				q			<=			16'h86B3;
		end
		32'h0000D762: begin
				q			<=			16'h00B6;
		end
		32'h0000D764: begin
				q			<=			16'hA683;
		end
		32'h0000D766: begin
				q			<=			16'hFE06;
		end
		32'h0000D768: begin
				q			<=			16'h0813;
		end
		32'h0000D76A: begin
				q			<=			16'h0200;
		end
		32'h0000D76C: begin
				q			<=			16'h0833;
		end
		32'h0000D76E: begin
				q			<=			16'h40E8;
		end
		32'h0000D770: begin
				q			<=			16'h96B3;
		end
		32'h0000D772: begin
				q			<=			16'h0106;
		end
		32'h0000D774: begin
				q			<=			16'h6633;
		end
		32'h0000D776: begin
				q			<=			16'h00D6;
		end
		32'h0000D778: begin
				q			<=			16'h0693;
		end
		32'h0000D77A: begin
				q			<=			16'h0030;
		end
		32'h0000D77C: begin
				q			<=			16'h0E13;
		end
		32'h0000D77E: begin
				q			<=			16'h0000;
		end
		32'h0000D780: begin
				q			<=			16'h86B3;
		end
		32'h0000D782: begin
				q			<=			16'h40F6;
		end
		32'h0000D784: begin
				q			<=			16'h4463;
		end
		32'h0000D786: begin
				q			<=			16'h02DE;
		end
		32'h0000D788: begin
				q			<=			16'h0593;
		end
		32'h0000D78A: begin
				q			<=			16'h0040;
		end
		32'h0000D78C: begin
				q			<=			16'h87B3;
		end
		32'h0000D78E: begin
				q			<=			16'h40F5;
		end
		32'h0000D790: begin
				q			<=			16'h9693;
		end
		32'h0000D792: begin
				q			<=			16'h0026;
		end
		32'h0000D794: begin
				q			<=			16'h0593;
		end
		32'h0000D796: begin
				q			<=			16'h0401;
		end
		32'h0000D798: begin
				q			<=			16'h86B3;
		end
		32'h0000D79A: begin
				q			<=			16'h00D5;
		end
		32'h0000D79C: begin
				q			<=			16'h2583;
		end
		32'h0000D79E: begin
				q			<=			16'h02C1;
		end
		32'h0000D7A0: begin
				q			<=			16'hD733;
		end
		32'h0000D7A2: begin
				q			<=			16'h00E5;
		end
		32'h0000D7A4: begin
				q			<=			16'hA023;
		end
		32'h0000D7A6: begin
				q			<=			16'hFEE6;
		end
		32'h0000D7A8: begin
				q			<=			16'hF06F;
		end
		32'h0000D7AA: begin
				q			<=			16'hF05F;
		end
		32'h0000D7AC: begin
				q			<=			16'h0EB3;
		end
		32'h0000D7AE: begin
				q			<=			16'h00B3;
		end
		32'h0000D7B0: begin
				q			<=			16'hA503;
		end
		32'h0000D7B2: begin
				q			<=			16'h000E;
		end
		32'h0000D7B4: begin
				q			<=			16'hAE83;
		end
		32'h0000D7B6: begin
				q			<=			16'h004E;
		end
		32'h0000D7B8: begin
				q			<=			16'h0E13;
		end
		32'h0000D7BA: begin
				q			<=			16'h001E;
		end
		32'h0000D7BC: begin
				q			<=			16'h5533;
		end
		32'h0000D7BE: begin
				q			<=			16'h00E5;
		end
		32'h0000D7C0: begin
				q			<=			16'h9EB3;
		end
		32'h0000D7C2: begin
				q			<=			16'h010E;
		end
		32'h0000D7C4: begin
				q			<=			16'h6533;
		end
		32'h0000D7C6: begin
				q			<=			16'h01D5;
		end
		32'h0000D7C8: begin
				q			<=			16'h2023;
		end
		32'h0000D7CA: begin
				q			<=			16'h00A3;
		end
		32'h0000D7CC: begin
				q			<=			16'h0313;
		end
		32'h0000D7CE: begin
				q			<=			16'h0043;
		end
		32'h0000D7D0: begin
				q			<=			16'hF06F;
		end
		32'h0000D7D2: begin
				q			<=			16'hFB5F;
		end
		32'h0000D7D4: begin
				q			<=			16'h9713;
		end
		32'h0000D7D6: begin
				q			<=			16'h0027;
		end
		32'h0000D7D8: begin
				q			<=			16'h8733;
		end
		32'h0000D7DA: begin
				q			<=			16'h00E8;
		end
		32'h0000D7DC: begin
				q			<=			16'h2023;
		end
		32'h0000D7DE: begin
				q			<=			16'h0007;
		end
		32'h0000D7E0: begin
				q			<=			16'h8793;
		end
		32'h0000D7E2: begin
				q			<=			16'h0017;
		end
		32'h0000D7E4: begin
				q			<=			16'hF06F;
		end
		32'h0000D7E6: begin
				q			<=			16'hECDF;
		end
		32'h0000D7E8: begin
				q			<=			16'h0063;
		end
		32'h0000D7EA: begin
				q			<=			16'h3E07;
		end
		32'h0000D7EC: begin
				q			<=			16'h1663;
		end
		32'h0000D7EE: begin
				q			<=			16'h2404;
		end
		32'h0000D7F0: begin
				q			<=			16'h2883;
		end
		32'h0000D7F2: begin
				q			<=			16'h0141;
		end
		32'h0000D7F4: begin
				q			<=			16'h2503;
		end
		32'h0000D7F6: begin
				q			<=			16'h0181;
		end
		32'h0000D7F8: begin
				q			<=			16'h2E03;
		end
		32'h0000D7FA: begin
				q			<=			16'h01C1;
		end
		32'h0000D7FC: begin
				q			<=			16'hE333;
		end
		32'h0000D7FE: begin
				q			<=			16'h00A8;
		end
		32'h0000D800: begin
				q			<=			16'h6333;
		end
		32'h0000D802: begin
				q			<=			16'h01C3;
		end
		32'h0000D804: begin
				q			<=			16'h6333;
		end
		32'h0000D806: begin
				q			<=			16'h00D3;
		end
		32'h0000D808: begin
				q			<=			16'h1E63;
		end
		32'h0000D80A: begin
				q			<=			16'h1803;
		end
		32'h0000D80C: begin
				q			<=			16'h2823;
		end
		32'h0000D80E: begin
				q			<=			16'h02F1;
		end
		32'h0000D810: begin
				q			<=			16'h2783;
		end
		32'h0000D812: begin
				q			<=			16'h0241;
		end
		32'h0000D814: begin
				q			<=			16'h0413;
		end
		32'h0000D816: begin
				q			<=			16'h0006;
		end
		32'h0000D818: begin
				q			<=			16'h2A23;
		end
		32'h0000D81A: begin
				q			<=			16'h02F1;
		end
		32'h0000D81C: begin
				q			<=			16'h2783;
		end
		32'h0000D81E: begin
				q			<=			16'h0281;
		end
		32'h0000D820: begin
				q			<=			16'h2C23;
		end
		32'h0000D822: begin
				q			<=			16'h02F1;
		end
		32'h0000D824: begin
				q			<=			16'h2783;
		end
		32'h0000D826: begin
				q			<=			16'h02C1;
		end
		32'h0000D828: begin
				q			<=			16'h2E23;
		end
		32'h0000D82A: begin
				q			<=			16'h02F1;
		end
		32'h0000D82C: begin
				q			<=			16'h2783;
		end
		32'h0000D82E: begin
				q			<=			16'h0301;
		end
		32'h0000D830: begin
				q			<=			16'hF713;
		end
		32'h0000D832: begin
				q			<=			16'h0077;
		end
		32'h0000D834: begin
				q			<=			16'h0463;
		end
		32'h0000D836: begin
				q			<=			16'h0407;
		end
		32'h0000D838: begin
				q			<=			16'hF713;
		end
		32'h0000D83A: begin
				q			<=			16'h00F7;
		end
		32'h0000D83C: begin
				q			<=			16'h0693;
		end
		32'h0000D83E: begin
				q			<=			16'h0040;
		end
		32'h0000D840: begin
				q			<=			16'h0E63;
		end
		32'h0000D842: begin
				q			<=			16'h02D7;
		end
		32'h0000D844: begin
				q			<=			16'h2703;
		end
		32'h0000D846: begin
				q			<=			16'h0341;
		end
		32'h0000D848: begin
				q			<=			16'h8793;
		end
		32'h0000D84A: begin
				q			<=			16'h0047;
		end
		32'h0000D84C: begin
				q			<=			16'h2823;
		end
		32'h0000D84E: begin
				q			<=			16'h02F1;
		end
		32'h0000D850: begin
				q			<=			16'hB793;
		end
		32'h0000D852: begin
				q			<=			16'h0047;
		end
		32'h0000D854: begin
				q			<=			16'h8733;
		end
		32'h0000D856: begin
				q			<=			16'h00E7;
		end
		32'h0000D858: begin
				q			<=			16'h37B3;
		end
		32'h0000D85A: begin
				q			<=			16'h00F7;
		end
		32'h0000D85C: begin
				q			<=			16'h2A23;
		end
		32'h0000D85E: begin
				q			<=			16'h02E1;
		end
		32'h0000D860: begin
				q			<=			16'h2703;
		end
		32'h0000D862: begin
				q			<=			16'h0381;
		end
		32'h0000D864: begin
				q			<=			16'h8733;
		end
		32'h0000D866: begin
				q			<=			16'h00E7;
		end
		32'h0000D868: begin
				q			<=			16'h2C23;
		end
		32'h0000D86A: begin
				q			<=			16'h02E1;
		end
		32'h0000D86C: begin
				q			<=			16'h3733;
		end
		32'h0000D86E: begin
				q			<=			16'h00F7;
		end
		32'h0000D870: begin
				q			<=			16'h2783;
		end
		32'h0000D872: begin
				q			<=			16'h03C1;
		end
		32'h0000D874: begin
				q			<=			16'h0733;
		end
		32'h0000D876: begin
				q			<=			16'h00F7;
		end
		32'h0000D878: begin
				q			<=			16'h2E23;
		end
		32'h0000D87A: begin
				q			<=			16'h02E1;
		end
		32'h0000D87C: begin
				q			<=			16'h2783;
		end
		32'h0000D87E: begin
				q			<=			16'h03C1;
		end
		32'h0000D880: begin
				q			<=			16'h9713;
		end
		32'h0000D882: begin
				q			<=			16'h00C7;
		end
		32'h0000D884: begin
				q			<=			16'h5263;
		end
		32'h0000D886: begin
				q			<=			16'h0207;
		end
		32'h0000D888: begin
				q			<=			16'h8737;
		end
		32'h0000D88A: begin
				q			<=			16'h0000;
		end
		32'h0000D88C: begin
				q			<=			16'h0413;
		end
		32'h0000D88E: begin
				q			<=			16'h0014;
		end
		32'h0000D890: begin
				q			<=			16'h0713;
		end
		32'h0000D892: begin
				q			<=			16'hFFF7;
		end
		32'h0000D894: begin
				q			<=			16'h08E3;
		end
		32'h0000D896: begin
				q			<=			16'h7AE4;
		end
		32'h0000D898: begin
				q			<=			16'h0737;
		end
		32'h0000D89A: begin
				q			<=			16'hFFF8;
		end
		32'h0000D89C: begin
				q			<=			16'h0713;
		end
		32'h0000D89E: begin
				q			<=			16'hFFF7;
		end
		32'h0000D8A0: begin
				q			<=			16'hF7B3;
		end
		32'h0000D8A2: begin
				q			<=			16'h00E7;
		end
		32'h0000D8A4: begin
				q			<=			16'h2E23;
		end
		32'h0000D8A6: begin
				q			<=			16'h02F1;
		end
		32'h0000D8A8: begin
				q			<=			16'h0793;
		end
		32'h0000D8AA: begin
				q			<=			16'h0301;
		end
		32'h0000D8AC: begin
				q			<=			16'h0693;
		end
		32'h0000D8AE: begin
				q			<=			16'h0000;
		end
		32'h0000D8B0: begin
				q			<=			16'h0593;
		end
		32'h0000D8B2: begin
				q			<=			16'h0030;
		end
		32'h0000D8B4: begin
				q			<=			16'hA703;
		end
		32'h0000D8B6: begin
				q			<=			16'h0007;
		end
		32'h0000D8B8: begin
				q			<=			16'hA603;
		end
		32'h0000D8BA: begin
				q			<=			16'h0047;
		end
		32'h0000D8BC: begin
				q			<=			16'h8693;
		end
		32'h0000D8BE: begin
				q			<=			16'h0016;
		end
		32'h0000D8C0: begin
				q			<=			16'h5713;
		end
		32'h0000D8C2: begin
				q			<=			16'h0037;
		end
		32'h0000D8C4: begin
				q			<=			16'h1613;
		end
		32'h0000D8C6: begin
				q			<=			16'h01D6;
		end
		32'h0000D8C8: begin
				q			<=			16'h6733;
		end
		32'h0000D8CA: begin
				q			<=			16'h00C7;
		end
		32'h0000D8CC: begin
				q			<=			16'hA023;
		end
		32'h0000D8CE: begin
				q			<=			16'h00E7;
		end
		32'h0000D8D0: begin
				q			<=			16'h8793;
		end
		32'h0000D8D2: begin
				q			<=			16'h0047;
		end
		32'h0000D8D4: begin
				q			<=			16'h90E3;
		end
		32'h0000D8D6: begin
				q			<=			16'hFEB6;
		end
		32'h0000D8D8: begin
				q			<=			16'h2783;
		end
		32'h0000D8DA: begin
				q			<=			16'h03C1;
		end
		32'h0000D8DC: begin
				q			<=			16'h86B7;
		end
		32'h0000D8DE: begin
				q			<=			16'h0000;
		end
		32'h0000D8E0: begin
				q			<=			16'hD713;
		end
		32'h0000D8E2: begin
				q			<=			16'h0037;
		end
		32'h0000D8E4: begin
				q			<=			16'h2E23;
		end
		32'h0000D8E6: begin
				q			<=			16'h02E1;
		end
		32'h0000D8E8: begin
				q			<=			16'h8793;
		end
		32'h0000D8EA: begin
				q			<=			16'hFFF6;
		end
		32'h0000D8EC: begin
				q			<=			16'h1A63;
		end
		32'h0000D8EE: begin
				q			<=			16'h02F4;
		end
		32'h0000D8F0: begin
				q			<=			16'h2603;
		end
		32'h0000D8F2: begin
				q			<=			16'h0341;
		end
		32'h0000D8F4: begin
				q			<=			16'h2783;
		end
		32'h0000D8F6: begin
				q			<=			16'h0301;
		end
		32'h0000D8F8: begin
				q			<=			16'hE7B3;
		end
		32'h0000D8FA: begin
				q			<=			16'h00C7;
		end
		32'h0000D8FC: begin
				q			<=			16'h2603;
		end
		32'h0000D8FE: begin
				q			<=			16'h0381;
		end
		32'h0000D900: begin
				q			<=			16'hE7B3;
		end
		32'h0000D902: begin
				q			<=			16'h00C7;
		end
		32'h0000D904: begin
				q			<=			16'hE7B3;
		end
		32'h0000D906: begin
				q			<=			16'h00E7;
		end
		32'h0000D908: begin
				q			<=			16'h8C63;
		end
		32'h0000D90A: begin
				q			<=			16'h0007;
		end
		32'h0000D90C: begin
				q			<=			16'h2E23;
		end
		32'h0000D90E: begin
				q			<=			16'h02D1;
		end
		32'h0000D910: begin
				q			<=			16'h2C23;
		end
		32'h0000D912: begin
				q			<=			16'h0201;
		end
		32'h0000D914: begin
				q			<=			16'h2A23;
		end
		32'h0000D916: begin
				q			<=			16'h0201;
		end
		32'h0000D918: begin
				q			<=			16'h2823;
		end
		32'h0000D91A: begin
				q			<=			16'h0201;
		end
		32'h0000D91C: begin
				q			<=			16'h0913;
		end
		32'h0000D91E: begin
				q			<=			16'h0000;
		end
		32'h0000D920: begin
				q			<=			16'h8537;
		end
		32'h0000D922: begin
				q			<=			16'h0000;
		end
		32'h0000D924: begin
				q			<=			16'h2783;
		end
		32'h0000D926: begin
				q			<=			16'h03C1;
		end
		32'h0000D928: begin
				q			<=			16'h0513;
		end
		32'h0000D92A: begin
				q			<=			16'hFFF5;
		end
		32'h0000D92C: begin
				q			<=			16'h7533;
		end
		32'h0000D92E: begin
				q			<=			16'h00A4;
		end
		32'h0000D930: begin
				q			<=			16'h5403;
		end
		32'h0000D932: begin
				q			<=			16'h00E1;
		end
		32'h0000D934: begin
				q			<=			16'h1623;
		end
		32'h0000D936: begin
				q			<=			16'h00F1;
		end
		32'h0000D938: begin
				q			<=			16'h87B7;
		end
		32'h0000D93A: begin
				q			<=			16'hFFFF;
		end
		32'h0000D93C: begin
				q			<=			16'h7433;
		end
		32'h0000D93E: begin
				q			<=			16'h00F4;
		end
		32'h0000D940: begin
				q			<=			16'h6433;
		end
		32'h0000D942: begin
				q			<=			16'h00A4;
		end
		32'h0000D944: begin
				q			<=			16'h5793;
		end
		32'h0000D946: begin
				q			<=			16'h0084;
		end
		32'h0000D948: begin
				q			<=			16'h1713;
		end
		32'h0000D94A: begin
				q			<=			16'h0079;
		end
		32'h0000D94C: begin
				q			<=			16'hF913;
		end
		32'h0000D94E: begin
				q			<=			16'h07F7;
		end
		32'h0000D950: begin
				q			<=			16'h2783;
		end
		32'h0000D952: begin
				q			<=			16'h0301;
		end
		32'h0000D954: begin
				q			<=			16'h1723;
		end
		32'h0000D956: begin
				q			<=			16'h0081;
		end
		32'h0000D958: begin
				q			<=			16'h6933;
		end
		32'h0000D95A: begin
				q			<=			16'h00E9;
		end
		32'h0000D95C: begin
				q			<=			16'hA023;
		end
		32'h0000D95E: begin
				q			<=			16'h00F4;
		end
		32'h0000D960: begin
				q			<=			16'h2783;
		end
		32'h0000D962: begin
				q			<=			16'h0341;
		end
		32'h0000D964: begin
				q			<=			16'h07A3;
		end
		32'h0000D966: begin
				q			<=			16'h0121;
		end
		32'h0000D968: begin
				q			<=			16'h2083;
		end
		32'h0000D96A: begin
				q			<=			16'h05C1;
		end
		32'h0000D96C: begin
				q			<=			16'hA223;
		end
		32'h0000D96E: begin
				q			<=			16'h00F4;
		end
		32'h0000D970: begin
				q			<=			16'h2783;
		end
		32'h0000D972: begin
				q			<=			16'h0381;
		end
		32'h0000D974: begin
				q			<=			16'h2403;
		end
		32'h0000D976: begin
				q			<=			16'h0581;
		end
		32'h0000D978: begin
				q			<=			16'h8513;
		end
		32'h0000D97A: begin
				q			<=			16'h0004;
		end
		32'h0000D97C: begin
				q			<=			16'hA423;
		end
		32'h0000D97E: begin
				q			<=			16'h00F4;
		end
		32'h0000D980: begin
				q			<=			16'h2783;
		end
		32'h0000D982: begin
				q			<=			16'h00C1;
		end
		32'h0000D984: begin
				q			<=			16'h2903;
		end
		32'h0000D986: begin
				q			<=			16'h0501;
		end
		32'h0000D988: begin
				q			<=			16'h2983;
		end
		32'h0000D98A: begin
				q			<=			16'h04C1;
		end
		32'h0000D98C: begin
				q			<=			16'hA623;
		end
		32'h0000D98E: begin
				q			<=			16'h00F4;
		end
		32'h0000D990: begin
				q			<=			16'h2A03;
		end
		32'h0000D992: begin
				q			<=			16'h0481;
		end
		32'h0000D994: begin
				q			<=			16'h2483;
		end
		32'h0000D996: begin
				q			<=			16'h0541;
		end
		32'h0000D998: begin
				q			<=			16'h2A83;
		end
		32'h0000D99A: begin
				q			<=			16'h0441;
		end
		32'h0000D99C: begin
				q			<=			16'h0113;
		end
		32'h0000D99E: begin
				q			<=			16'h0601;
		end
		32'h0000D9A0: begin
				q			<=			16'h8067;
		end
		32'h0000D9A2: begin
				q			<=			16'h0000;
		end
		32'h0000D9A4: begin
				q			<=			16'h0313;
		end
		32'h0000D9A6: begin
				q			<=			16'hFFF0;
		end
		32'h0000D9A8: begin
				q			<=			16'h1063;
		end
		32'h0000D9AA: begin
				q			<=			16'h0667;
		end
		32'h0000D9AC: begin
				q			<=			16'h2583;
		end
		32'h0000D9AE: begin
				q			<=			16'h0241;
		end
		32'h0000D9B0: begin
				q			<=			16'h86B3;
		end
		32'h0000D9B2: begin
				q			<=			16'h00F6;
		end
		32'h0000D9B4: begin
				q			<=			16'hB7B3;
		end
		32'h0000D9B6: begin
				q			<=			16'h00F6;
		end
		32'h0000D9B8: begin
				q			<=			16'h8833;
		end
		32'h0000D9BA: begin
				q			<=			16'h00B8;
		end
		32'h0000D9BC: begin
				q			<=			16'h0733;
		end
		32'h0000D9BE: begin
				q			<=			16'h00F8;
		end
		32'h0000D9C0: begin
				q			<=			16'h37B3;
		end
		32'h0000D9C2: begin
				q			<=			16'h00F7;
		end
		32'h0000D9C4: begin
				q			<=			16'h2A23;
		end
		32'h0000D9C6: begin
				q			<=			16'h02E1;
		end
		32'h0000D9C8: begin
				q			<=			16'h2703;
		end
		32'h0000D9CA: begin
				q			<=			16'h0281;
		end
		32'h0000D9CC: begin
				q			<=			16'h35B3;
		end
		32'h0000D9CE: begin
				q			<=			16'h00B8;
		end
		32'h0000D9D0: begin
				q			<=			16'hE7B3;
		end
		32'h0000D9D2: begin
				q			<=			16'h00F5;
		end
		32'h0000D9D4: begin
				q			<=			16'h2823;
		end
		32'h0000D9D6: begin
				q			<=			16'h02D1;
		end
		32'h0000D9D8: begin
				q			<=			16'h06B3;
		end
		32'h0000D9DA: begin
				q			<=			16'h00E5;
		end
		32'h0000D9DC: begin
				q			<=			16'h85B3;
		end
		32'h0000D9DE: begin
				q			<=			16'h00F6;
		end
		32'h0000D9E0: begin
				q			<=			16'hB7B3;
		end
		32'h0000D9E2: begin
				q			<=			16'h00F5;
		end
		32'h0000D9E4: begin
				q			<=			16'hB733;
		end
		32'h0000D9E6: begin
				q			<=			16'h00E6;
		end
		32'h0000D9E8: begin
				q			<=			16'h6733;
		end
		32'h0000D9EA: begin
				q			<=			16'h00F7;
		end
		32'h0000D9EC: begin
				q			<=			16'h2783;
		end
		32'h0000D9EE: begin
				q			<=			16'h02C1;
		end
		32'h0000D9F0: begin
				q			<=			16'h2C23;
		end
		32'h0000D9F2: begin
				q			<=			16'h02B1;
		end
		32'h0000D9F4: begin
				q			<=			16'h0E33;
		end
		32'h0000D9F6: begin
				q			<=			16'h00FE;
		end
		32'h0000D9F8: begin
				q			<=			16'h0733;
		end
		32'h0000D9FA: begin
				q			<=			16'h01C7;
		end
		32'h0000D9FC: begin
				q			<=			16'h2E23;
		end
		32'h0000D9FE: begin
				q			<=			16'h02E1;
		end
		32'h0000DA00: begin
				q			<=			16'h0413;
		end
		32'h0000DA02: begin
				q			<=			16'h0006;
		end
		32'h0000DA04: begin
				q			<=			16'hF06F;
		end
		32'h0000DA06: begin
				q			<=			16'hB85F;
		end
		32'h0000DA08: begin
				q			<=			16'h86B7;
		end
		32'h0000DA0A: begin
				q			<=			16'h0000;
		end
		32'h0000DA0C: begin
				q			<=			16'h8693;
		end
		32'h0000DA0E: begin
				q			<=			16'hFFF6;
		end
		32'h0000DA10: begin
				q			<=			16'h0EE3;
		end
		32'h0000DA12: begin
				q			<=			16'hDED6;
		end
		32'h0000DA14: begin
				q			<=			16'h4713;
		end
		32'h0000DA16: begin
				q			<=			16'hFFF7;
		end
		32'h0000DA18: begin
				q			<=			16'h0793;
		end
		32'h0000DA1A: begin
				q			<=			16'h0740;
		end
		32'h0000DA1C: begin
				q			<=			16'hD263;
		end
		32'h0000DA1E: begin
				q			<=			16'h04E7;
		end
		32'h0000DA20: begin
				q			<=			16'h0793;
		end
		32'h0000DA22: begin
				q			<=			16'h0010;
		end
		32'h0000DA24: begin
				q			<=			16'h2E23;
		end
		32'h0000DA26: begin
				q			<=			16'h0001;
		end
		32'h0000DA28: begin
				q			<=			16'h2C23;
		end
		32'h0000DA2A: begin
				q			<=			16'h0001;
		end
		32'h0000DA2C: begin
				q			<=			16'h2A23;
		end
		32'h0000DA2E: begin
				q			<=			16'h0001;
		end
		32'h0000DA30: begin
				q			<=			16'h2823;
		end
		32'h0000DA32: begin
				q			<=			16'h00F1;
		end
		32'h0000DA34: begin
				q			<=			16'h006F;
		end
		32'h0000DA36: begin
				q			<=			16'h0740;
		end
		32'h0000DA38: begin
				q			<=			16'h86B7;
		end
		32'h0000DA3A: begin
				q			<=			16'h0000;
		end
		32'h0000DA3C: begin
				q			<=			16'h8693;
		end
		32'h0000DA3E: begin
				q			<=			16'hFFF6;
		end
		32'h0000DA40: begin
				q			<=			16'h06E3;
		end
		32'h0000DA42: begin
				q			<=			16'hDCD6;
		end
		32'h0000DA44: begin
				q			<=			16'h2783;
		end
		32'h0000DA46: begin
				q			<=			16'h01C1;
		end
		32'h0000DA48: begin
				q			<=			16'h06B7;
		end
		32'h0000DA4A: begin
				q			<=			16'h0008;
		end
		32'h0000DA4C: begin
				q			<=			16'hE7B3;
		end
		32'h0000DA4E: begin
				q			<=			16'h00D7;
		end
		32'h0000DA50: begin
				q			<=			16'h2E23;
		end
		32'h0000DA52: begin
				q			<=			16'h00F1;
		end
		32'h0000DA54: begin
				q			<=			16'h0793;
		end
		32'h0000DA56: begin
				q			<=			16'hF8C0;
		end
		32'h0000DA58: begin
				q			<=			16'h44E3;
		end
		32'h0000DA5A: begin
				q			<=			16'hFCF7;
		end
		32'h0000DA5C: begin
				q			<=			16'h0733;
		end
		32'h0000DA5E: begin
				q			<=			16'h40E0;
		end
		32'h0000DA60: begin
				q			<=			16'h5693;
		end
		32'h0000DA62: begin
				q			<=			16'h4057;
		end
		32'h0000DA64: begin
				q			<=			16'h0513;
		end
		32'h0000DA66: begin
				q			<=			16'h0000;
		end
		32'h0000DA68: begin
				q			<=			16'h7713;
		end
		32'h0000DA6A: begin
				q			<=			16'h01F7;
		end
		32'h0000DA6C: begin
				q			<=			16'h0793;
		end
		32'h0000DA6E: begin
				q			<=			16'h0000;
		end
		32'h0000DA70: begin
				q			<=			16'h9893;
		end
		32'h0000DA72: begin
				q			<=			16'h0027;
		end
		32'h0000DA74: begin
				q			<=			16'h9E63;
		end
		32'h0000DA76: begin
				q			<=			16'h08D7;
		end
		32'h0000DA78: begin
				q			<=			16'h1263;
		end
		32'h0000DA7A: begin
				q			<=			16'h0C07;
		end
		32'h0000DA7C: begin
				q			<=			16'h0693;
		end
		32'h0000DA7E: begin
				q			<=			16'h0030;
		end
		32'h0000DA80: begin
				q			<=			16'h86B3;
		end
		32'h0000DA82: begin
				q			<=			16'h40F6;
		end
		32'h0000DA84: begin
				q			<=			16'hD063;
		end
		32'h0000DA86: begin
				q			<=			16'h0AE6;
		end
		32'h0000DA88: begin
				q			<=			16'h0713;
		end
		32'h0000DA8A: begin
				q			<=			16'h0040;
		end
		32'h0000DA8C: begin
				q			<=			16'h07B3;
		end
		32'h0000DA8E: begin
				q			<=			16'h40F7;
		end
		32'h0000DA90: begin
				q			<=			16'h0693;
		end
		32'h0000DA92: begin
				q			<=			16'h0040;
		end
		32'h0000DA94: begin
				q			<=			16'h9063;
		end
		32'h0000DA96: begin
				q			<=			16'h12D7;
		end
		32'h0000DA98: begin
				q			<=			16'h2783;
		end
		32'h0000DA9A: begin
				q			<=			16'h0101;
		end
		32'h0000DA9C: begin
				q			<=			16'h3533;
		end
		32'h0000DA9E: begin
				q			<=			16'h00A0;
		end
		32'h0000DAA0: begin
				q			<=			16'hE533;
		end
		32'h0000DAA2: begin
				q			<=			16'h00A7;
		end
		32'h0000DAA4: begin
				q			<=			16'h2823;
		end
		32'h0000DAA6: begin
				q			<=			16'h00A1;
		end
		32'h0000DAA8: begin
				q			<=			16'h2683;
		end
		32'h0000DAAA: begin
				q			<=			16'h0201;
		end
		32'h0000DAAC: begin
				q			<=			16'h2783;
		end
		32'h0000DAAE: begin
				q			<=			16'h0101;
		end
		32'h0000DAB0: begin
				q			<=			16'h2703;
		end
		32'h0000DAB2: begin
				q			<=			16'h0241;
		end
		32'h0000DAB4: begin
				q			<=			16'h2503;
		end
		32'h0000DAB6: begin
				q			<=			16'h0181;
		end
		32'h0000DAB8: begin
				q			<=			16'h87B3;
		end
		32'h0000DABA: begin
				q			<=			16'h00F6;
		end
		32'h0000DABC: begin
				q			<=			16'hB6B3;
		end
		32'h0000DABE: begin
				q			<=			16'h00D7;
		end
		32'h0000DAC0: begin
				q			<=			16'h2823;
		end
		32'h0000DAC2: begin
				q			<=			16'h02F1;
		end
		32'h0000DAC4: begin
				q			<=			16'h2783;
		end
		32'h0000DAC6: begin
				q			<=			16'h0141;
		end
		32'h0000DAC8: begin
				q			<=			16'h2803;
		end
		32'h0000DACA: begin
				q			<=			16'h01C1;
		end
		32'h0000DACC: begin
				q			<=			16'h07B3;
		end
		32'h0000DACE: begin
				q			<=			16'h00F7;
		end
		32'h0000DAD0: begin
				q			<=			16'h85B3;
		end
		32'h0000DAD2: begin
				q			<=			16'h00D7;
		end
		32'h0000DAD4: begin
				q			<=			16'hB733;
		end
		32'h0000DAD6: begin
				q			<=			16'h00E7;
		end
		32'h0000DAD8: begin
				q			<=			16'hB7B3;
		end
		32'h0000DADA: begin
				q			<=			16'h00D5;
		end
		32'h0000DADC: begin
				q			<=			16'h67B3;
		end
		32'h0000DADE: begin
				q			<=			16'h00F7;
		end
		32'h0000DAE0: begin
				q			<=			16'h2703;
		end
		32'h0000DAE2: begin
				q			<=			16'h0281;
		end
		32'h0000DAE4: begin
				q			<=			16'h2683;
		end
		32'h0000DAE6: begin
				q			<=			16'h02C1;
		end
		32'h0000DAE8: begin
				q			<=			16'h2A23;
		end
		32'h0000DAEA: begin
				q			<=			16'h02B1;
		end
		32'h0000DAEC: begin
				q			<=			16'h0533;
		end
		32'h0000DAEE: begin
				q			<=			16'h00A7;
		end
		32'h0000DAF0: begin
				q			<=			16'h05B3;
		end
		32'h0000DAF2: begin
				q			<=			16'h00F5;
		end
		32'h0000DAF4: begin
				q			<=			16'h3733;
		end
		32'h0000DAF6: begin
				q			<=			16'h00E5;
		end
		32'h0000DAF8: begin
				q			<=			16'hB7B3;
		end
		32'h0000DAFA: begin
				q			<=			16'h00F5;
		end
		32'h0000DAFC: begin
				q			<=			16'h86B3;
		end
		32'h0000DAFE: begin
				q			<=			16'h0106;
		end
		32'h0000DB00: begin
				q			<=			16'h6733;
		end
		32'h0000DB02: begin
				q			<=			16'h00F7;
		end
		32'h0000DB04: begin
				q			<=			16'h2C23;
		end
		32'h0000DB06: begin
				q			<=			16'h02B1;
		end
		32'h0000DB08: begin
				q			<=			16'h8733;
		end
		32'h0000DB0A: begin
				q			<=			16'h00E6;
		end
		32'h0000DB0C: begin
				q			<=			16'hF06F;
		end
		32'h0000DB0E: begin
				q			<=			16'hEF1F;
		end
		32'h0000DB10: begin
				q			<=			16'h08B3;
		end
		32'h0000DB12: begin
				q			<=			16'h0118;
		end
		32'h0000DB14: begin
				q			<=			16'hA883;
		end
		32'h0000DB16: begin
				q			<=			16'h0008;
		end
		32'h0000DB18: begin
				q			<=			16'h8793;
		end
		32'h0000DB1A: begin
				q			<=			16'h0017;
		end
		32'h0000DB1C: begin
				q			<=			16'h6533;
		end
		32'h0000DB1E: begin
				q			<=			16'h0115;
		end
		32'h0000DB20: begin
				q			<=			16'hF06F;
		end
		32'h0000DB22: begin
				q			<=			16'hF51F;
		end
		32'h0000DB24: begin
				q			<=			16'h8333;
		end
		32'h0000DB26: begin
				q			<=			16'h0115;
		end
		32'h0000DB28: begin
				q			<=			16'h2303;
		end
		32'h0000DB2A: begin
				q			<=			16'h0003;
		end
		32'h0000DB2C: begin
				q			<=			16'h0713;
		end
		32'h0000DB2E: begin
				q			<=			16'h0017;
		end
		32'h0000DB30: begin
				q			<=			16'h8593;
		end
		32'h0000DB32: begin
				q			<=			16'h0045;
		end
		32'h0000DB34: begin
				q			<=			16'hAE23;
		end
		32'h0000DB36: begin
				q			<=			16'hFE65;
		end
		32'h0000DB38: begin
				q			<=			16'hF06F;
		end
		32'h0000DB3A: begin
				q			<=			16'hF4DF;
		end
		32'h0000DB3C: begin
				q			<=			16'h0693;
		end
		32'h0000DB3E: begin
				q			<=			16'h0401;
		end
		32'h0000DB40: begin
				q			<=			16'h86B3;
		end
		32'h0000DB42: begin
				q			<=			16'h0116;
		end
		32'h0000DB44: begin
				q			<=			16'hA683;
		end
		32'h0000DB46: begin
				q			<=			16'hFD06;
		end
		32'h0000DB48: begin
				q			<=			16'h0E13;
		end
		32'h0000DB4A: begin
				q			<=			16'h0200;
		end
		32'h0000DB4C: begin
				q			<=			16'h0E33;
		end
		32'h0000DB4E: begin
				q			<=			16'h40EE;
		end
		32'h0000DB50: begin
				q			<=			16'h96B3;
		end
		32'h0000DB52: begin
				q			<=			16'h01C6;
		end
		32'h0000DB54: begin
				q			<=			16'h6533;
		end
		32'h0000DB56: begin
				q			<=			16'h00D5;
		end
		32'h0000DB58: begin
				q			<=			16'h0693;
		end
		32'h0000DB5A: begin
				q			<=			16'h0030;
		end
		32'h0000DB5C: begin
				q			<=			16'h0E93;
		end
		32'h0000DB5E: begin
				q			<=			16'h0000;
		end
		32'h0000DB60: begin
				q			<=			16'h86B3;
		end
		32'h0000DB62: begin
				q			<=			16'h40F6;
		end
		32'h0000DB64: begin
				q			<=			16'hC463;
		end
		32'h0000DB66: begin
				q			<=			16'h02DE;
		end
		32'h0000DB68: begin
				q			<=			16'h0593;
		end
		32'h0000DB6A: begin
				q			<=			16'h0040;
		end
		32'h0000DB6C: begin
				q			<=			16'h87B3;
		end
		32'h0000DB6E: begin
				q			<=			16'h40F5;
		end
		32'h0000DB70: begin
				q			<=			16'h9693;
		end
		32'h0000DB72: begin
				q			<=			16'h0026;
		end
		32'h0000DB74: begin
				q			<=			16'h0593;
		end
		32'h0000DB76: begin
				q			<=			16'h0401;
		end
		32'h0000DB78: begin
				q			<=			16'h86B3;
		end
		32'h0000DB7A: begin
				q			<=			16'h00D5;
		end
		32'h0000DB7C: begin
				q			<=			16'h2583;
		end
		32'h0000DB7E: begin
				q			<=			16'h01C1;
		end
		32'h0000DB80: begin
				q			<=			16'hD733;
		end
		32'h0000DB82: begin
				q			<=			16'h00E5;
		end
		32'h0000DB84: begin
				q			<=			16'hA823;
		end
		32'h0000DB86: begin
				q			<=			16'hFCE6;
		end
		32'h0000DB88: begin
				q			<=			16'hF06F;
		end
		32'h0000DB8A: begin
				q			<=			16'hF09F;
		end
		32'h0000DB8C: begin
				q			<=			16'h8F33;
		end
		32'h0000DB8E: begin
				q			<=			16'h0115;
		end
		32'h0000DB90: begin
				q			<=			16'h2303;
		end
		32'h0000DB92: begin
				q			<=			16'h000F;
		end
		32'h0000DB94: begin
				q			<=			16'h2F03;
		end
		32'h0000DB96: begin
				q			<=			16'h004F;
		end
		32'h0000DB98: begin
				q			<=			16'h8E93;
		end
		32'h0000DB9A: begin
				q			<=			16'h001E;
		end
		32'h0000DB9C: begin
				q			<=			16'h5333;
		end
		32'h0000DB9E: begin
				q			<=			16'h00E3;
		end
		32'h0000DBA0: begin
				q			<=			16'h1F33;
		end
		32'h0000DBA2: begin
				q			<=			16'h01CF;
		end
		32'h0000DBA4: begin
				q			<=			16'h6333;
		end
		32'h0000DBA6: begin
				q			<=			16'h01E3;
		end
		32'h0000DBA8: begin
				q			<=			16'hA023;
		end
		32'h0000DBAA: begin
				q			<=			16'h0065;
		end
		32'h0000DBAC: begin
				q			<=			16'h8593;
		end
		32'h0000DBAE: begin
				q			<=			16'h0045;
		end
		32'h0000DBB0: begin
				q			<=			16'hF06F;
		end
		32'h0000DBB2: begin
				q			<=			16'hFB5F;
		end
		32'h0000DBB4: begin
				q			<=			16'h9713;
		end
		32'h0000DBB6: begin
				q			<=			16'h0027;
		end
		32'h0000DBB8: begin
				q			<=			16'h0733;
		end
		32'h0000DBBA: begin
				q			<=			16'h00E8;
		end
		32'h0000DBBC: begin
				q			<=			16'h2023;
		end
		32'h0000DBBE: begin
				q			<=			16'h0007;
		end
		32'h0000DBC0: begin
				q			<=			16'h8793;
		end
		32'h0000DBC2: begin
				q			<=			16'h0017;
		end
		32'h0000DBC4: begin
				q			<=			16'hF06F;
		end
		32'h0000DBC6: begin
				q			<=			16'hED1F;
		end
		32'h0000DBC8: begin
				q			<=			16'h8F37;
		end
		32'h0000DBCA: begin
				q			<=			16'h0000;
		end
		32'h0000DBCC: begin
				q			<=			16'h0593;
		end
		32'h0000DBCE: begin
				q			<=			16'h0014;
		end
		32'h0000DBD0: begin
				q			<=			16'h0E93;
		end
		32'h0000DBD2: begin
				q			<=			16'hFFFF;
		end
		32'h0000DBD4: begin
				q			<=			16'hF2B3;
		end
		32'h0000DBD6: begin
				q			<=			16'h01D5;
		end
		32'h0000DBD8: begin
				q			<=			16'h0F93;
		end
		32'h0000DBDA: begin
				q			<=			16'h0010;
		end
		32'h0000DBDC: begin
				q			<=			16'h2603;
		end
		32'h0000DBDE: begin
				q			<=			16'h0241;
		end
		32'h0000DBE0: begin
				q			<=			16'h2703;
		end
		32'h0000DBE2: begin
				q			<=			16'h0281;
		end
		32'h0000DBE4: begin
				q			<=			16'h2503;
		end
		32'h0000DBE6: begin
				q			<=			16'h02C1;
		end
		32'h0000DBE8: begin
				q			<=			16'h2E03;
		end
		32'h0000DBEA: begin
				q			<=			16'h0141;
		end
		32'h0000DBEC: begin
				q			<=			16'h2883;
		end
		32'h0000DBEE: begin
				q			<=			16'h0181;
		end
		32'h0000DBF0: begin
				q			<=			16'h2303;
		end
		32'h0000DBF2: begin
				q			<=			16'h01C1;
		end
		32'h0000DBF4: begin
				q			<=			16'h0813;
		end
		32'h0000DBF6: begin
				q			<=			16'h0301;
		end
		32'h0000DBF8: begin
				q			<=			16'hC663;
		end
		32'h0000DBFA: begin
				q			<=			16'h145F;
		end
		32'h0000DBFC: begin
				q			<=			16'h65B3;
		end
		32'h0000DBFE: begin
				q			<=			16'h011E;
		end
		32'h0000DC00: begin
				q			<=			16'hE5B3;
		end
		32'h0000DC02: begin
				q			<=			16'h0065;
		end
		32'h0000DC04: begin
				q			<=			16'hE5B3;
		end
		32'h0000DC06: begin
				q			<=			16'h00D5;
		end
		32'h0000DC08: begin
				q			<=			16'h1663;
		end
		32'h0000DC0A: begin
				q			<=			16'h0A04;
		end
		32'h0000DC0C: begin
				q			<=			16'h9C63;
		end
		32'h0000DC0E: begin
				q			<=			16'h0005;
		end
		32'h0000DC10: begin
				q			<=			16'h2823;
		end
		32'h0000DC12: begin
				q			<=			16'h02F1;
		end
		32'h0000DC14: begin
				q			<=			16'h2A23;
		end
		32'h0000DC16: begin
				q			<=			16'h02C1;
		end
		32'h0000DC18: begin
				q			<=			16'h2C23;
		end
		32'h0000DC1A: begin
				q			<=			16'h02E1;
		end
		32'h0000DC1C: begin
				q			<=			16'h2E23;
		end
		32'h0000DC1E: begin
				q			<=			16'h02A1;
		end
		32'h0000DC20: begin
				q			<=			16'hF06F;
		end
		32'h0000DC22: begin
				q			<=			16'hC0DF;
		end
		32'h0000DC24: begin
				q			<=			16'h65B3;
		end
		32'h0000DC26: begin
				q			<=			16'h00E6;
		end
		32'h0000DC28: begin
				q			<=			16'hE5B3;
		end
		32'h0000DC2A: begin
				q			<=			16'h00A5;
		end
		32'h0000DC2C: begin
				q			<=			16'hE5B3;
		end
		32'h0000DC2E: begin
				q			<=			16'h00F5;
		end
		32'h0000DC30: begin
				q			<=			16'h9C63;
		end
		32'h0000DC32: begin
				q			<=			16'h0005;
		end
		32'h0000DC34: begin
				q			<=			16'h2823;
		end
		32'h0000DC36: begin
				q			<=			16'h02D1;
		end
		32'h0000DC38: begin
				q			<=			16'h2A23;
		end
		32'h0000DC3A: begin
				q			<=			16'h03C1;
		end
		32'h0000DC3C: begin
				q			<=			16'h2C23;
		end
		32'h0000DC3E: begin
				q			<=			16'h0311;
		end
		32'h0000DC40: begin
				q			<=			16'h2E23;
		end
		32'h0000DC42: begin
				q			<=			16'h0261;
		end
		32'h0000DC44: begin
				q			<=			16'hF06F;
		end
		32'h0000DC46: begin
				q			<=			16'hBE9F;
		end
		32'h0000DC48: begin
				q			<=			16'h87B3;
		end
		32'h0000DC4A: begin
				q			<=			16'h00F6;
		end
		32'h0000DC4C: begin
				q			<=			16'h0633;
		end
		32'h0000DC4E: begin
				q			<=			16'h01C6;
		end
		32'h0000DC50: begin
				q			<=			16'h2823;
		end
		32'h0000DC52: begin
				q			<=			16'h02F1;
		end
		32'h0000DC54: begin
				q			<=			16'hB7B3;
		end
		32'h0000DC56: begin
				q			<=			16'h00D7;
		end
		32'h0000DC58: begin
				q			<=			16'h06B3;
		end
		32'h0000DC5A: begin
				q			<=			16'h00F6;
		end
		32'h0000DC5C: begin
				q			<=			16'h2A23;
		end
		32'h0000DC5E: begin
				q			<=			16'h02D1;
		end
		32'h0000DC60: begin
				q			<=			16'h3633;
		end
		32'h0000DC62: begin
				q			<=			16'h01C6;
		end
		32'h0000DC64: begin
				q			<=			16'hB6B3;
		end
		32'h0000DC66: begin
				q			<=			16'h00F6;
		end
		32'h0000DC68: begin
				q			<=			16'h66B3;
		end
		32'h0000DC6A: begin
				q			<=			16'h00D6;
		end
		32'h0000DC6C: begin
				q			<=			16'h05B3;
		end
		32'h0000DC6E: begin
				q			<=			16'h0117;
		end
		32'h0000DC70: begin
				q			<=			16'h87B3;
		end
		32'h0000DC72: begin
				q			<=			16'h00D5;
		end
		32'h0000DC74: begin
				q			<=			16'hB733;
		end
		32'h0000DC76: begin
				q			<=			16'h0115;
		end
		32'h0000DC78: begin
				q			<=			16'hB6B3;
		end
		32'h0000DC7A: begin
				q			<=			16'h00D7;
		end
		32'h0000DC7C: begin
				q			<=			16'h66B3;
		end
		32'h0000DC7E: begin
				q			<=			16'h00D7;
		end
		32'h0000DC80: begin
				q			<=			16'h0733;
		end
		32'h0000DC82: begin
				q			<=			16'h0065;
		end
		32'h0000DC84: begin
				q			<=			16'h8733;
		end
		32'h0000DC86: begin
				q			<=			16'h00E6;
		end
		32'h0000DC88: begin
				q			<=			16'h2C23;
		end
		32'h0000DC8A: begin
				q			<=			16'h02F1;
		end
		32'h0000DC8C: begin
				q			<=			16'h1793;
		end
		32'h0000DC8E: begin
				q			<=			16'h00C7;
		end
		32'h0000DC90: begin
				q			<=			16'hC663;
		end
		32'h0000DC92: begin
				q			<=			16'h0007;
		end
		32'h0000DC94: begin
				q			<=			16'h2E23;
		end
		32'h0000DC96: begin
				q			<=			16'h02E1;
		end
		32'h0000DC98: begin
				q			<=			16'hF06F;
		end
		32'h0000DC9A: begin
				q			<=			16'hB95F;
		end
		32'h0000DC9C: begin
				q			<=			16'h06B7;
		end
		32'h0000DC9E: begin
				q			<=			16'hFFF8;
		end
		32'h0000DCA0: begin
				q			<=			16'h8693;
		end
		32'h0000DCA2: begin
				q			<=			16'hFFF6;
		end
		32'h0000DCA4: begin
				q			<=			16'h7733;
		end
		32'h0000DCA6: begin
				q			<=			16'h00D7;
		end
		32'h0000DCA8: begin
				q			<=			16'h2E23;
		end
		32'h0000DCAA: begin
				q			<=			16'h02E1;
		end
		32'h0000DCAC: begin
				q			<=			16'h0413;
		end
		32'h0000DCAE: begin
				q			<=			16'h0010;
		end
		32'h0000DCB0: begin
				q			<=			16'hF06F;
		end
		32'h0000DCB2: begin
				q			<=			16'hB7DF;
		end
		32'h0000DCB4: begin
				q			<=			16'h9E63;
		end
		32'h0000DCB6: begin
				q			<=			16'h0005;
		end
		32'h0000DCB8: begin
				q			<=			16'h2823;
		end
		32'h0000DCBA: begin
				q			<=			16'h02F1;
		end
		32'h0000DCBC: begin
				q			<=			16'h2A23;
		end
		32'h0000DCBE: begin
				q			<=			16'h02C1;
		end
		32'h0000DCC0: begin
				q			<=			16'h2C23;
		end
		32'h0000DCC2: begin
				q			<=			16'h02E1;
		end
		32'h0000DCC4: begin
				q			<=			16'h2E23;
		end
		32'h0000DCC6: begin
				q			<=			16'h02A1;
		end
		32'h0000DCC8: begin
				q			<=			16'h8413;
		end
		32'h0000DCCA: begin
				q			<=			16'h000E;
		end
		32'h0000DCCC: begin
				q			<=			16'hF06F;
		end
		32'h0000DCCE: begin
				q			<=			16'hB61F;
		end
		32'h0000DCD0: begin
				q			<=			16'h6733;
		end
		32'h0000DCD2: begin
				q			<=			16'h00E6;
		end
		32'h0000DCD4: begin
				q			<=			16'h6733;
		end
		32'h0000DCD6: begin
				q			<=			16'h00A7;
		end
		32'h0000DCD8: begin
				q			<=			16'h67B3;
		end
		32'h0000DCDA: begin
				q			<=			16'h00F7;
		end
		32'h0000DCDC: begin
				q			<=			16'h9C63;
		end
		32'h0000DCDE: begin
				q			<=			16'h0007;
		end
		32'h0000DCE0: begin
				q			<=			16'h2823;
		end
		32'h0000DCE2: begin
				q			<=			16'h02D1;
		end
		32'h0000DCE4: begin
				q			<=			16'h2A23;
		end
		32'h0000DCE6: begin
				q			<=			16'h03C1;
		end
		32'h0000DCE8: begin
				q			<=			16'h2C23;
		end
		32'h0000DCEA: begin
				q			<=			16'h0311;
		end
		32'h0000DCEC: begin
				q			<=			16'h2E23;
		end
		32'h0000DCEE: begin
				q			<=			16'h0261;
		end
		32'h0000DCF0: begin
				q			<=			16'hF06F;
		end
		32'h0000DCF2: begin
				q			<=			16'hFD9F;
		end
		32'h0000DCF4: begin
				q			<=			16'h2E23;
		end
		32'h0000DCF6: begin
				q			<=			16'h03E1;
		end
		32'h0000DCF8: begin
				q			<=			16'h2C23;
		end
		32'h0000DCFA: begin
				q			<=			16'h0201;
		end
		32'h0000DCFC: begin
				q			<=			16'h2A23;
		end
		32'h0000DCFE: begin
				q			<=			16'h0201;
		end
		32'h0000DD00: begin
				q			<=			16'h2823;
		end
		32'h0000DD02: begin
				q			<=			16'h0201;
		end
		32'h0000DD04: begin
				q			<=			16'h0793;
		end
		32'h0000DD06: begin
				q			<=			16'h03C1;
		end
		32'h0000DD08: begin
				q			<=			16'hA703;
		end
		32'h0000DD0A: begin
				q			<=			16'h0007;
		end
		32'h0000DD0C: begin
				q			<=			16'hA683;
		end
		32'h0000DD0E: begin
				q			<=			16'hFFC7;
		end
		32'h0000DD10: begin
				q			<=			16'h8793;
		end
		32'h0000DD12: begin
				q			<=			16'hFFC7;
		end
		32'h0000DD14: begin
				q			<=			16'h1713;
		end
		32'h0000DD16: begin
				q			<=			16'h0037;
		end
		32'h0000DD18: begin
				q			<=			16'hD693;
		end
		32'h0000DD1A: begin
				q			<=			16'h01D6;
		end
		32'h0000DD1C: begin
				q			<=			16'h6733;
		end
		32'h0000DD1E: begin
				q			<=			16'h00D7;
		end
		32'h0000DD20: begin
				q			<=			16'hA223;
		end
		32'h0000DD22: begin
				q			<=			16'h00E7;
		end
		32'h0000DD24: begin
				q			<=			16'h12E3;
		end
		32'h0000DD26: begin
				q			<=			16'hFEF8;
		end
		32'h0000DD28: begin
				q			<=			16'h2783;
		end
		32'h0000DD2A: begin
				q			<=			16'h0301;
		end
		32'h0000DD2C: begin
				q			<=			16'h8437;
		end
		32'h0000DD2E: begin
				q			<=			16'h0000;
		end
		32'h0000DD30: begin
				q			<=			16'h0413;
		end
		32'h0000DD32: begin
				q			<=			16'hFFF4;
		end
		32'h0000DD34: begin
				q			<=			16'h9793;
		end
		32'h0000DD36: begin
				q			<=			16'h0037;
		end
		32'h0000DD38: begin
				q			<=			16'h2823;
		end
		32'h0000DD3A: begin
				q			<=			16'h02F1;
		end
		32'h0000DD3C: begin
				q			<=			16'h0913;
		end
		32'h0000DD3E: begin
				q			<=			16'h0000;
		end
		32'h0000DD40: begin
				q			<=			16'hF06F;
		end
		32'h0000DD42: begin
				q			<=			16'hAEDF;
		end
		32'h0000DD44: begin
				q			<=			16'h87B3;
		end
		32'h0000DD46: begin
				q			<=			16'h00F6;
		end
		32'h0000DD48: begin
				q			<=			16'h0633;
		end
		32'h0000DD4A: begin
				q			<=			16'h01C6;
		end
		32'h0000DD4C: begin
				q			<=			16'h2823;
		end
		32'h0000DD4E: begin
				q			<=			16'h02F1;
		end
		32'h0000DD50: begin
				q			<=			16'hB7B3;
		end
		32'h0000DD52: begin
				q			<=			16'h00D7;
		end
		32'h0000DD54: begin
				q			<=			16'h06B3;
		end
		32'h0000DD56: begin
				q			<=			16'h00F6;
		end
		32'h0000DD58: begin
				q			<=			16'h2A23;
		end
		32'h0000DD5A: begin
				q			<=			16'h02D1;
		end
		32'h0000DD5C: begin
				q			<=			16'h3633;
		end
		32'h0000DD5E: begin
				q			<=			16'h01C6;
		end
		32'h0000DD60: begin
				q			<=			16'hB6B3;
		end
		32'h0000DD62: begin
				q			<=			16'h00F6;
		end
		32'h0000DD64: begin
				q			<=			16'h66B3;
		end
		32'h0000DD66: begin
				q			<=			16'h00D6;
		end
		32'h0000DD68: begin
				q			<=			16'h0733;
		end
		32'h0000DD6A: begin
				q			<=			16'h0117;
		end
		32'h0000DD6C: begin
				q			<=			16'h0633;
		end
		32'h0000DD6E: begin
				q			<=			16'h00D7;
		end
		32'h0000DD70: begin
				q			<=			16'h36B3;
		end
		32'h0000DD72: begin
				q			<=			16'h00D6;
		end
		32'h0000DD74: begin
				q			<=			16'h3733;
		end
		32'h0000DD76: begin
				q			<=			16'h0117;
		end
		32'h0000DD78: begin
				q			<=			16'h66B3;
		end
		32'h0000DD7A: begin
				q			<=			16'h00D7;
		end
		32'h0000DD7C: begin
				q			<=			16'h0733;
		end
		32'h0000DD7E: begin
				q			<=			16'h0065;
		end
		32'h0000DD80: begin
				q			<=			16'h8733;
		end
		32'h0000DD82: begin
				q			<=			16'h00E6;
		end
		32'h0000DD84: begin
				q			<=			16'h2C23;
		end
		32'h0000DD86: begin
				q			<=			16'h02C1;
		end
		32'h0000DD88: begin
				q			<=			16'h2E23;
		end
		32'h0000DD8A: begin
				q			<=			16'h02E1;
		end
		32'h0000DD8C: begin
				q			<=			16'h0793;
		end
		32'h0000DD8E: begin
				q			<=			16'h0008;
		end
		32'h0000DD90: begin
				q			<=			16'h0693;
		end
		32'h0000DD92: begin
				q			<=			16'h0000;
		end
		32'h0000DD94: begin
				q			<=			16'h0513;
		end
		32'h0000DD96: begin
				q			<=			16'h0030;
		end
		32'h0000DD98: begin
				q			<=			16'hA703;
		end
		32'h0000DD9A: begin
				q			<=			16'h0007;
		end
		32'h0000DD9C: begin
				q			<=			16'hA603;
		end
		32'h0000DD9E: begin
				q			<=			16'h0047;
		end
		32'h0000DDA0: begin
				q			<=			16'h8693;
		end
		32'h0000DDA2: begin
				q			<=			16'h0016;
		end
		32'h0000DDA4: begin
				q			<=			16'h5713;
		end
		32'h0000DDA6: begin
				q			<=			16'h0017;
		end
		32'h0000DDA8: begin
				q			<=			16'h1613;
		end
		32'h0000DDAA: begin
				q			<=			16'h01F6;
		end
		32'h0000DDAC: begin
				q			<=			16'h6733;
		end
		32'h0000DDAE: begin
				q			<=			16'h00C7;
		end
		32'h0000DDB0: begin
				q			<=			16'hA023;
		end
		32'h0000DDB2: begin
				q			<=			16'h00E7;
		end
		32'h0000DDB4: begin
				q			<=			16'h8793;
		end
		32'h0000DDB6: begin
				q			<=			16'h0047;
		end
		32'h0000DDB8: begin
				q			<=			16'h90E3;
		end
		32'h0000DDBA: begin
				q			<=			16'hFEA6;
		end
		32'h0000DDBC: begin
				q			<=			16'h2783;
		end
		32'h0000DDBE: begin
				q			<=			16'h03C1;
		end
		32'h0000DDC0: begin
				q			<=			16'h8413;
		end
		32'h0000DDC2: begin
				q			<=			16'h0005;
		end
		32'h0000DDC4: begin
				q			<=			16'hD793;
		end
		32'h0000DDC6: begin
				q			<=			16'h0017;
		end
		32'h0000DDC8: begin
				q			<=			16'h2E23;
		end
		32'h0000DDCA: begin
				q			<=			16'h02F1;
		end
		32'h0000DDCC: begin
				q			<=			16'h87B7;
		end
		32'h0000DDCE: begin
				q			<=			16'h0000;
		end
		32'h0000DDD0: begin
				q			<=			16'h8793;
		end
		32'h0000DDD2: begin
				q			<=			16'hFFF7;
		end
		32'h0000DDD4: begin
				q			<=			16'h1CE3;
		end
		32'h0000DDD6: begin
				q			<=			16'hA4F4;
		end
		32'h0000DDD8: begin
				q			<=			16'h2E23;
		end
		32'h0000DDDA: begin
				q			<=			16'h0201;
		end
		32'h0000DDDC: begin
				q			<=			16'h2C23;
		end
		32'h0000DDDE: begin
				q			<=			16'h0201;
		end
		32'h0000DDE0: begin
				q			<=			16'h2A23;
		end
		32'h0000DDE2: begin
				q			<=			16'h0201;
		end
		32'h0000DDE4: begin
				q			<=			16'h2823;
		end
		32'h0000DDE6: begin
				q			<=			16'h0201;
		end
		32'h0000DDE8: begin
				q			<=			16'hF06F;
		end
		32'h0000DDEA: begin
				q			<=			16'hA45F;
		end
		32'h0000DDEC: begin
				q			<=			16'h5463;
		end
		32'h0000DDEE: begin
				q			<=			16'h28E0;
		end
		32'h0000DDF0: begin
				q			<=			16'h1063;
		end
		32'h0000DDF2: begin
				q			<=			16'h0E06;
		end
		32'h0000DDF4: begin
				q			<=			16'h2503;
		end
		32'h0000DDF6: begin
				q			<=			16'h0241;
		end
		32'h0000DDF8: begin
				q			<=			16'h2583;
		end
		32'h0000DDFA: begin
				q			<=			16'h0281;
		end
		32'h0000DDFC: begin
				q			<=			16'h2E03;
		end
		32'h0000DDFE: begin
				q			<=			16'h02C1;
		end
		32'h0000DE00: begin
				q			<=			16'h6833;
		end
		32'h0000DE02: begin
				q			<=			16'h00B5;
		end
		32'h0000DE04: begin
				q			<=			16'h6833;
		end
		32'h0000DE06: begin
				q			<=			16'h01C8;
		end
		32'h0000DE08: begin
				q			<=			16'h6833;
		end
		32'h0000DE0A: begin
				q			<=			16'h00F8;
		end
		32'h0000DE0C: begin
				q			<=			16'h0C63;
		end
		32'h0000DE0E: begin
				q			<=			16'hEE08;
		end
		32'h0000DE10: begin
				q			<=			16'h0613;
		end
		32'h0000DE12: begin
				q			<=			16'hFFF7;
		end
		32'h0000DE14: begin
				q			<=			16'h1863;
		end
		32'h0000DE16: begin
				q			<=			16'h0806;
		end
		32'h0000DE18: begin
				q			<=			16'h2883;
		end
		32'h0000DE1A: begin
				q			<=			16'h0141;
		end
		32'h0000DE1C: begin
				q			<=			16'h87B3;
		end
		32'h0000DE1E: begin
				q			<=			16'h40F6;
		end
		32'h0000DE20: begin
				q			<=			16'hB733;
		end
		32'h0000DE22: begin
				q			<=			16'h00F6;
		end
		32'h0000DE24: begin
				q			<=			16'h8833;
		end
		32'h0000DE26: begin
				q			<=			16'h40A8;
		end
		32'h0000DE28: begin
				q			<=			16'hB333;
		end
		32'h0000DE2A: begin
				q			<=			16'h0108;
		end
		32'h0000DE2C: begin
				q			<=			16'h0833;
		end
		32'h0000DE2E: begin
				q			<=			16'h40E8;
		end
		32'h0000DE30: begin
				q			<=			16'h2823;
		end
		32'h0000DE32: begin
				q			<=			16'h02F1;
		end
		32'h0000DE34: begin
				q			<=			16'h2A23;
		end
		32'h0000DE36: begin
				q			<=			16'h0301;
		end
		32'h0000DE38: begin
				q			<=			16'h0713;
		end
		32'h0000DE3A: begin
				q			<=			16'h0000;
		end
		32'h0000DE3C: begin
				q			<=			16'hF663;
		end
		32'h0000DE3E: begin
				q			<=			16'h00F6;
		end
		32'h0000DE40: begin
				q			<=			16'h0733;
		end
		32'h0000DE42: begin
				q			<=			16'h4115;
		end
		32'h0000DE44: begin
				q			<=			16'h3713;
		end
		32'h0000DE46: begin
				q			<=			16'h0017;
		end
		32'h0000DE48: begin
				q			<=			16'h2803;
		end
		32'h0000DE4A: begin
				q			<=			16'h0181;
		end
		32'h0000DE4C: begin
				q			<=			16'h6733;
		end
		32'h0000DE4E: begin
				q			<=			16'h0067;
		end
		32'h0000DE50: begin
				q			<=			16'h06B3;
		end
		32'h0000DE52: begin
				q			<=			16'h40B8;
		end
		32'h0000DE54: begin
				q			<=			16'h3533;
		end
		32'h0000DE56: begin
				q			<=			16'h00D8;
		end
		32'h0000DE58: begin
				q			<=			16'h86B3;
		end
		32'h0000DE5A: begin
				q			<=			16'h40E6;
		end
		32'h0000DE5C: begin
				q			<=			16'h2C23;
		end
		32'h0000DE5E: begin
				q			<=			16'h02D1;
		end
		32'h0000DE60: begin
				q			<=			16'h0663;
		end
		32'h0000DE62: begin
				q			<=			16'h0007;
		end
		32'h0000DE64: begin
				q			<=			16'h85B3;
		end
		32'h0000DE66: begin
				q			<=			16'h4105;
		end
		32'h0000DE68: begin
				q			<=			16'hB613;
		end
		32'h0000DE6A: begin
				q			<=			16'h0015;
		end
		32'h0000DE6C: begin
				q			<=			16'h2783;
		end
		32'h0000DE6E: begin
				q			<=			16'h01C1;
		end
		32'h0000DE70: begin
				q			<=			16'h6633;
		end
		32'h0000DE72: begin
				q			<=			16'h00A6;
		end
		32'h0000DE74: begin
				q			<=			16'h0413;
		end
		32'h0000DE76: begin
				q			<=			16'h0010;
		end
		32'h0000DE78: begin
				q			<=			16'h87B3;
		end
		32'h0000DE7A: begin
				q			<=			16'h41C7;
		end
		32'h0000DE7C: begin
				q			<=			16'h8633;
		end
		32'h0000DE7E: begin
				q			<=			16'h40C7;
		end
		32'h0000DE80: begin
				q			<=			16'h2E23;
		end
		32'h0000DE82: begin
				q			<=			16'h02C1;
		end
		32'h0000DE84: begin
				q			<=			16'h2783;
		end
		32'h0000DE86: begin
				q			<=			16'h03C1;
		end
		32'h0000DE88: begin
				q			<=			16'h9713;
		end
		32'h0000DE8A: begin
				q			<=			16'h00C7;
		end
		32'h0000DE8C: begin
				q			<=			16'h50E3;
		end
		32'h0000DE8E: begin
				q			<=			16'h9A07;
		end
		32'h0000DE90: begin
				q			<=			16'h0737;
		end
		32'h0000DE92: begin
				q			<=			16'h0008;
		end
		32'h0000DE94: begin
				q			<=			16'h0713;
		end
		32'h0000DE96: begin
				q			<=			16'hFFF7;
		end
		32'h0000DE98: begin
				q			<=			16'hF7B3;
		end
		32'h0000DE9A: begin
				q			<=			16'h00E7;
		end
		32'h0000DE9C: begin
				q			<=			16'h2E23;
		end
		32'h0000DE9E: begin
				q			<=			16'h02F1;
		end
		32'h0000DEA0: begin
				q			<=			16'h006F;
		end
		32'h0000DEA2: begin
				q			<=			16'h7340;
		end
		32'h0000DEA4: begin
				q			<=			16'h87B7;
		end
		32'h0000DEA6: begin
				q			<=			16'h0000;
		end
		32'h0000DEA8: begin
				q			<=			16'h8793;
		end
		32'h0000DEAA: begin
				q			<=			16'hFFF7;
		end
		32'h0000DEAC: begin
				q			<=			16'h0C63;
		end
		32'h0000DEAE: begin
				q			<=			16'hE4F7;
		end
		32'h0000DEB0: begin
				q			<=			16'h0793;
		end
		32'h0000DEB2: begin
				q			<=			16'h0740;
		end
		32'h0000DEB4: begin
				q			<=			16'hD263;
		end
		32'h0000DEB6: begin
				q			<=			16'h04C7;
		end
		32'h0000DEB8: begin
				q			<=			16'h0793;
		end
		32'h0000DEBA: begin
				q			<=			16'h0010;
		end
		32'h0000DEBC: begin
				q			<=			16'h2623;
		end
		32'h0000DEBE: begin
				q			<=			16'h0201;
		end
		32'h0000DEC0: begin
				q			<=			16'h2423;
		end
		32'h0000DEC2: begin
				q			<=			16'h0201;
		end
		32'h0000DEC4: begin
				q			<=			16'h2223;
		end
		32'h0000DEC6: begin
				q			<=			16'h0201;
		end
		32'h0000DEC8: begin
				q			<=			16'h2023;
		end
		32'h0000DECA: begin
				q			<=			16'h02F1;
		end
		32'h0000DECC: begin
				q			<=			16'h006F;
		end
		32'h0000DECE: begin
				q			<=			16'h0740;
		end
		32'h0000DED0: begin
				q			<=			16'h87B7;
		end
		32'h0000DED2: begin
				q			<=			16'h0000;
		end
		32'h0000DED4: begin
				q			<=			16'h8793;
		end
		32'h0000DED6: begin
				q			<=			16'hFFF7;
		end
		32'h0000DED8: begin
				q			<=			16'h0463;
		end
		32'h0000DEDA: begin
				q			<=			16'hF6F4;
		end
		32'h0000DEDC: begin
				q			<=			16'h2783;
		end
		32'h0000DEDE: begin
				q			<=			16'h02C1;
		end
		32'h0000DEE0: begin
				q			<=			16'h06B7;
		end
		32'h0000DEE2: begin
				q			<=			16'h0008;
		end
		32'h0000DEE4: begin
				q			<=			16'hE7B3;
		end
		32'h0000DEE6: begin
				q			<=			16'h00D7;
		end
		32'h0000DEE8: begin
				q			<=			16'h2623;
		end
		32'h0000DEEA: begin
				q			<=			16'h02F1;
		end
		32'h0000DEEC: begin
				q			<=			16'h0793;
		end
		32'h0000DEEE: begin
				q			<=			16'h0740;
		end
		32'h0000DEF0: begin
				q			<=			16'hC4E3;
		end
		32'h0000DEF2: begin
				q			<=			16'hFCE7;
		end
		32'h0000DEF4: begin
				q			<=			16'h0613;
		end
		32'h0000DEF6: begin
				q			<=			16'h0007;
		end
		32'h0000DEF8: begin
				q			<=			16'h5713;
		end
		32'h0000DEFA: begin
				q			<=			16'h4056;
		end
		32'h0000DEFC: begin
				q			<=			16'h0693;
		end
		32'h0000DEFE: begin
				q			<=			16'h0000;
		end
		32'h0000DF00: begin
				q			<=			16'h7613;
		end
		32'h0000DF02: begin
				q			<=			16'h01F6;
		end
		32'h0000DF04: begin
				q			<=			16'h0793;
		end
		32'h0000DF06: begin
				q			<=			16'h0000;
		end
		32'h0000DF08: begin
				q			<=			16'h9593;
		end
		32'h0000DF0A: begin
				q			<=			16'h0027;
		end
		32'h0000DF0C: begin
				q			<=			16'h9863;
		end
		32'h0000DF0E: begin
				q			<=			16'h0AE7;
		end
		32'h0000DF10: begin
				q			<=			16'h1C63;
		end
		32'h0000DF12: begin
				q			<=			16'h0C06;
		end
		32'h0000DF14: begin
				q			<=			16'h0713;
		end
		32'h0000DF16: begin
				q			<=			16'h0030;
		end
		32'h0000DF18: begin
				q			<=			16'h0733;
		end
		32'h0000DF1A: begin
				q			<=			16'h40F7;
		end
		32'h0000DF1C: begin
				q			<=			16'h5A63;
		end
		32'h0000DF1E: begin
				q			<=			16'h0AC7;
		end
		32'h0000DF20: begin
				q			<=			16'h0713;
		end
		32'h0000DF22: begin
				q			<=			16'h0040;
		end
		32'h0000DF24: begin
				q			<=			16'h07B3;
		end
		32'h0000DF26: begin
				q			<=			16'h40F7;
		end
		32'h0000DF28: begin
				q			<=			16'h0613;
		end
		32'h0000DF2A: begin
				q			<=			16'h0040;
		end
		32'h0000DF2C: begin
				q			<=			16'h9A63;
		end
		32'h0000DF2E: begin
				q			<=			16'h12C7;
		end
		32'h0000DF30: begin
				q			<=			16'h2783;
		end
		32'h0000DF32: begin
				q			<=			16'h0201;
		end
		32'h0000DF34: begin
				q			<=			16'h36B3;
		end
		32'h0000DF36: begin
				q			<=			16'h00D0;
		end
		32'h0000DF38: begin
				q			<=			16'hE6B3;
		end
		32'h0000DF3A: begin
				q			<=			16'h00D7;
		end
		32'h0000DF3C: begin
				q			<=			16'h2023;
		end
		32'h0000DF3E: begin
				q			<=			16'h02D1;
		end
		32'h0000DF40: begin
				q			<=			16'h2683;
		end
		32'h0000DF42: begin
				q			<=			16'h0141;
		end
		32'h0000DF44: begin
				q			<=			16'h2583;
		end
		32'h0000DF46: begin
				q			<=			16'h0101;
		end
		32'h0000DF48: begin
				q			<=			16'h2703;
		end
		32'h0000DF4A: begin
				q			<=			16'h0201;
		end
		32'h0000DF4C: begin
				q			<=			16'h2783;
		end
		32'h0000DF4E: begin
				q			<=			16'h0241;
		end
		32'h0000DF50: begin
				q			<=			16'h8733;
		end
		32'h0000DF52: begin
				q			<=			16'h40E5;
		end
		32'h0000DF54: begin
				q			<=			16'h87B3;
		end
		32'h0000DF56: begin
				q			<=			16'h40F6;
		end
		32'h0000DF58: begin
				q			<=			16'hB633;
		end
		32'h0000DF5A: begin
				q			<=			16'h00F6;
		end
		32'h0000DF5C: begin
				q			<=			16'hB6B3;
		end
		32'h0000DF5E: begin
				q			<=			16'h00E5;
		end
		32'h0000DF60: begin
				q			<=			16'h86B3;
		end
		32'h0000DF62: begin
				q			<=			16'h40D7;
		end
		32'h0000DF64: begin
				q			<=			16'h2A23;
		end
		32'h0000DF66: begin
				q			<=			16'h02D1;
		end
		32'h0000DF68: begin
				q			<=			16'h2823;
		end
		32'h0000DF6A: begin
				q			<=			16'h02E1;
		end
		32'h0000DF6C: begin
				q			<=			16'h0693;
		end
		32'h0000DF6E: begin
				q			<=			16'h0000;
		end
		32'h0000DF70: begin
				q			<=			16'hF463;
		end
		32'h0000DF72: begin
				q			<=			16'h00E5;
		end
		32'h0000DF74: begin
				q			<=			16'hB693;
		end
		32'h0000DF76: begin
				q			<=			16'h0017;
		end
		32'h0000DF78: begin
				q			<=			16'hE6B3;
		end
		32'h0000DF7A: begin
				q			<=			16'h00C6;
		end
		32'h0000DF7C: begin
				q			<=			16'h2703;
		end
		32'h0000DF7E: begin
				q			<=			16'h0281;
		end
		32'h0000DF80: begin
				q			<=			16'h2603;
		end
		32'h0000DF82: begin
				q			<=			16'h0181;
		end
		32'h0000DF84: begin
				q			<=			16'h0733;
		end
		32'h0000DF86: begin
				q			<=			16'h40E6;
		end
		32'h0000DF88: begin
				q			<=			16'h07B3;
		end
		32'h0000DF8A: begin
				q			<=			16'h40D7;
		end
		32'h0000DF8C: begin
				q			<=			16'h2C23;
		end
		32'h0000DF8E: begin
				q			<=			16'h02F1;
		end
		32'h0000DF90: begin
				q			<=			16'h35B3;
		end
		32'h0000DF92: begin
				q			<=			16'h00E6;
		end
		32'h0000DF94: begin
				q			<=			16'h0613;
		end
		32'h0000DF96: begin
				q			<=			16'h0000;
		end
		32'h0000DF98: begin
				q			<=			16'h8463;
		end
		32'h0000DF9A: begin
				q			<=			16'h0006;
		end
		32'h0000DF9C: begin
				q			<=			16'h3613;
		end
		32'h0000DF9E: begin
				q			<=			16'h0017;
		end
		32'h0000DFA0: begin
				q			<=			16'h2783;
		end
		32'h0000DFA2: begin
				q			<=			16'h01C1;
		end
		32'h0000DFA4: begin
				q			<=			16'h2703;
		end
		32'h0000DFA6: begin
				q			<=			16'h02C1;
		end
		32'h0000DFA8: begin
				q			<=			16'h6633;
		end
		32'h0000DFAA: begin
				q			<=			16'h00B6;
		end
		32'h0000DFAC: begin
				q			<=			16'h87B3;
		end
		32'h0000DFAE: begin
				q			<=			16'h40E7;
		end
		32'h0000DFB0: begin
				q			<=			16'h87B3;
		end
		32'h0000DFB2: begin
				q			<=			16'h40C7;
		end
		32'h0000DFB4: begin
				q			<=			16'h2E23;
		end
		32'h0000DFB6: begin
				q			<=			16'h02F1;
		end
		32'h0000DFB8: begin
				q			<=			16'hF06F;
		end
		32'h0000DFBA: begin
				q			<=			16'hECDF;
		end
		32'h0000DFBC: begin
				q			<=			16'h85B3;
		end
		32'h0000DFBE: begin
				q			<=			16'h00B8;
		end
		32'h0000DFC0: begin
				q			<=			16'hA583;
		end
		32'h0000DFC2: begin
				q			<=			16'h0005;
		end
		32'h0000DFC4: begin
				q			<=			16'h8793;
		end
		32'h0000DFC6: begin
				q			<=			16'h0017;
		end
		32'h0000DFC8: begin
				q			<=			16'hE6B3;
		end
		32'h0000DFCA: begin
				q			<=			16'h00B6;
		end
		32'h0000DFCC: begin
				q			<=			16'hF06F;
		end
		32'h0000DFCE: begin
				q			<=			16'hF3DF;
		end
		32'h0000DFD0: begin
				q			<=			16'h0533;
		end
		32'h0000DFD2: begin
				q			<=			16'h00B3;
		end
		32'h0000DFD4: begin
				q			<=			16'h2503;
		end
		32'h0000DFD6: begin
				q			<=			16'h0005;
		end
		32'h0000DFD8: begin
				q			<=			16'h0613;
		end
		32'h0000DFDA: begin
				q			<=			16'h0016;
		end
		32'h0000DFDC: begin
				q			<=			16'h0313;
		end
		32'h0000DFDE: begin
				q			<=			16'h0043;
		end
		32'h0000DFE0: begin
				q			<=			16'h2E23;
		end
		32'h0000DFE2: begin
				q			<=			16'hFEA3;
		end
		32'h0000DFE4: begin
				q			<=			16'hF06F;
		end
		32'h0000DFE6: begin
				q			<=			16'hF39F;
		end
		32'h0000DFE8: begin
				q			<=			16'h0713;
		end
		32'h0000DFEA: begin
				q			<=			16'h0401;
		end
		32'h0000DFEC: begin
				q			<=			16'h0733;
		end
		32'h0000DFEE: begin
				q			<=			16'h00B7;
		end
		32'h0000DFF0: begin
				q			<=			16'h2703;
		end
		32'h0000DFF2: begin
				q			<=			16'hFE07;
		end
		32'h0000DFF4: begin
				q			<=			16'h0813;
		end
		32'h0000DFF6: begin
				q			<=			16'h0200;
		end
		32'h0000DFF8: begin
				q			<=			16'h0833;
		end
		32'h0000DFFA: begin
				q			<=			16'h40C8;
		end
		32'h0000DFFC: begin
				q			<=			16'h1733;
		end
		32'h0000DFFE: begin
				q			<=			16'h0107;
		end
		32'h0000E000: begin
				q			<=			16'hE6B3;
		end
		32'h0000E002: begin
				q			<=			16'h00E6;
		end
		32'h0000E004: begin
				q			<=			16'h0713;
		end
		32'h0000E006: begin
				q			<=			16'h0030;
		end
		32'h0000E008: begin
				q			<=			16'h0E13;
		end
		32'h0000E00A: begin
				q			<=			16'h0000;
		end
		32'h0000E00C: begin
				q			<=			16'h0733;
		end
		32'h0000E00E: begin
				q			<=			16'h40F7;
		end
		32'h0000E010: begin
				q			<=			16'h4463;
		end
		32'h0000E012: begin
				q			<=			16'h02EE;
		end
		32'h0000E014: begin
				q			<=			16'h0593;
		end
		32'h0000E016: begin
				q			<=			16'h0040;
		end
		32'h0000E018: begin
				q			<=			16'h87B3;
		end
		32'h0000E01A: begin
				q			<=			16'h40F5;
		end
		32'h0000E01C: begin
				q			<=			16'h1713;
		end
		32'h0000E01E: begin
				q			<=			16'h0027;
		end
		32'h0000E020: begin
				q			<=			16'h0593;
		end
		32'h0000E022: begin
				q			<=			16'h0401;
		end
		32'h0000E024: begin
				q			<=			16'h8733;
		end
		32'h0000E026: begin
				q			<=			16'h00E5;
		end
		32'h0000E028: begin
				q			<=			16'h2583;
		end
		32'h0000E02A: begin
				q			<=			16'h02C1;
		end
		32'h0000E02C: begin
				q			<=			16'hD633;
		end
		32'h0000E02E: begin
				q			<=			16'h00C5;
		end
		32'h0000E030: begin
				q			<=			16'h2023;
		end
		32'h0000E032: begin
				q			<=			16'hFEC7;
		end
		32'h0000E034: begin
				q			<=			16'hF06F;
		end
		32'h0000E036: begin
				q			<=			16'hEF5F;
		end
		32'h0000E038: begin
				q			<=			16'h0EB3;
		end
		32'h0000E03A: begin
				q			<=			16'h00B3;
		end
		32'h0000E03C: begin
				q			<=			16'hA503;
		end
		32'h0000E03E: begin
				q			<=			16'h000E;
		end
		32'h0000E040: begin
				q			<=			16'hAE83;
		end
		32'h0000E042: begin
				q			<=			16'h004E;
		end
		32'h0000E044: begin
				q			<=			16'h0E13;
		end
		32'h0000E046: begin
				q			<=			16'h001E;
		end
		32'h0000E048: begin
				q			<=			16'h5533;
		end
		32'h0000E04A: begin
				q			<=			16'h00C5;
		end
		32'h0000E04C: begin
				q			<=			16'h9EB3;
		end
		32'h0000E04E: begin
				q			<=			16'h010E;
		end
		32'h0000E050: begin
				q			<=			16'h6533;
		end
		32'h0000E052: begin
				q			<=			16'h01D5;
		end
		32'h0000E054: begin
				q			<=			16'h2023;
		end
		32'h0000E056: begin
				q			<=			16'h00A3;
		end
		32'h0000E058: begin
				q			<=			16'h0313;
		end
		32'h0000E05A: begin
				q			<=			16'h0043;
		end
		32'h0000E05C: begin
				q			<=			16'hF06F;
		end
		32'h0000E05E: begin
				q			<=			16'hFB5F;
		end
		32'h0000E060: begin
				q			<=			16'h9713;
		end
		32'h0000E062: begin
				q			<=			16'h0027;
		end
		32'h0000E064: begin
				q			<=			16'h8733;
		end
		32'h0000E066: begin
				q			<=			16'h00E8;
		end
		32'h0000E068: begin
				q			<=			16'h2023;
		end
		32'h0000E06A: begin
				q			<=			16'h0007;
		end
		32'h0000E06C: begin
				q			<=			16'h8793;
		end
		32'h0000E06E: begin
				q			<=			16'h0017;
		end
		32'h0000E070: begin
				q			<=			16'hF06F;
		end
		32'h0000E072: begin
				q			<=			16'hEBDF;
		end
		32'h0000E074: begin
				q			<=			16'h0E63;
		end
		32'h0000E076: begin
				q			<=			16'h2807;
		end
		32'h0000E078: begin
				q			<=			16'h1C63;
		end
		32'h0000E07A: begin
				q			<=			16'h0E04;
		end
		32'h0000E07C: begin
				q			<=			16'h2303;
		end
		32'h0000E07E: begin
				q			<=			16'h0141;
		end
		32'h0000E080: begin
				q			<=			16'h2883;
		end
		32'h0000E082: begin
				q			<=			16'h0181;
		end
		32'h0000E084: begin
				q			<=			16'h2E83;
		end
		32'h0000E086: begin
				q			<=			16'h01C1;
		end
		32'h0000E088: begin
				q			<=			16'h6E33;
		end
		32'h0000E08A: begin
				q			<=			16'h0113;
		end
		32'h0000E08C: begin
				q			<=			16'h6E33;
		end
		32'h0000E08E: begin
				q			<=			16'h01DE;
		end
		32'h0000E090: begin
				q			<=			16'h6E33;
		end
		32'h0000E092: begin
				q			<=			16'h00DE;
		end
		32'h0000E094: begin
				q			<=			16'h1663;
		end
		32'h0000E096: begin
				q			<=			16'h020E;
		end
		32'h0000E098: begin
				q			<=			16'h2823;
		end
		32'h0000E09A: begin
				q			<=			16'h02F1;
		end
		32'h0000E09C: begin
				q			<=			16'h2783;
		end
		32'h0000E09E: begin
				q			<=			16'h0241;
		end
		32'h0000E0A0: begin
				q			<=			16'h0413;
		end
		32'h0000E0A2: begin
				q			<=			16'h0006;
		end
		32'h0000E0A4: begin
				q			<=			16'h2A23;
		end
		32'h0000E0A6: begin
				q			<=			16'h02F1;
		end
		32'h0000E0A8: begin
				q			<=			16'h2783;
		end
		32'h0000E0AA: begin
				q			<=			16'h0281;
		end
		32'h0000E0AC: begin
				q			<=			16'h2C23;
		end
		32'h0000E0AE: begin
				q			<=			16'h02F1;
		end
		32'h0000E0B0: begin
				q			<=			16'h2783;
		end
		32'h0000E0B2: begin
				q			<=			16'h02C1;
		end
		32'h0000E0B4: begin
				q			<=			16'h2E23;
		end
		32'h0000E0B6: begin
				q			<=			16'h02F1;
		end
		32'h0000E0B8: begin
				q			<=			16'h0913;
		end
		32'h0000E0BA: begin
				q			<=			16'h0005;
		end
		32'h0000E0BC: begin
				q			<=			16'hF06F;
		end
		32'h0000E0BE: begin
				q			<=			16'hF70F;
		end
		32'h0000E0C0: begin
				q			<=			16'h0E13;
		end
		32'h0000E0C2: begin
				q			<=			16'hFFF0;
		end
		32'h0000E0C4: begin
				q			<=			16'h1E63;
		end
		32'h0000E0C6: begin
				q			<=			16'h07C7;
		end
		32'h0000E0C8: begin
				q			<=			16'h2803;
		end
		32'h0000E0CA: begin
				q			<=			16'h0241;
		end
		32'h0000E0CC: begin
				q			<=			16'h86B3;
		end
		32'h0000E0CE: begin
				q			<=			16'h40D7;
		end
		32'h0000E0D0: begin
				q			<=			16'hB733;
		end
		32'h0000E0D2: begin
				q			<=			16'h00D7;
		end
		32'h0000E0D4: begin
				q			<=			16'h05B3;
		end
		32'h0000E0D6: begin
				q			<=			16'h4068;
		end
		32'h0000E0D8: begin
				q			<=			16'h3E33;
		end
		32'h0000E0DA: begin
				q			<=			16'h00B8;
		end
		32'h0000E0DC: begin
				q			<=			16'h85B3;
		end
		32'h0000E0DE: begin
				q			<=			16'h40E5;
		end
		32'h0000E0E0: begin
				q			<=			16'h2823;
		end
		32'h0000E0E2: begin
				q			<=			16'h02D1;
		end
		32'h0000E0E4: begin
				q			<=			16'h2A23;
		end
		32'h0000E0E6: begin
				q			<=			16'h02B1;
		end
		32'h0000E0E8: begin
				q			<=			16'h0713;
		end
		32'h0000E0EA: begin
				q			<=			16'h0000;
		end
		32'h0000E0EC: begin
				q			<=			16'hF663;
		end
		32'h0000E0EE: begin
				q			<=			16'h00D7;
		end
		32'h0000E0F0: begin
				q			<=			16'h0733;
		end
		32'h0000E0F2: begin
				q			<=			16'h4103;
		end
		32'h0000E0F4: begin
				q			<=			16'h3713;
		end
		32'h0000E0F6: begin
				q			<=			16'h0017;
		end
		32'h0000E0F8: begin
				q			<=			16'h2803;
		end
		32'h0000E0FA: begin
				q			<=			16'h0281;
		end
		32'h0000E0FC: begin
				q			<=			16'h6733;
		end
		32'h0000E0FE: begin
				q			<=			16'h01C7;
		end
		32'h0000E100: begin
				q			<=			16'h0693;
		end
		32'h0000E102: begin
				q			<=			16'h0000;
		end
		32'h0000E104: begin
				q			<=			16'h05B3;
		end
		32'h0000E106: begin
				q			<=			16'h4118;
		end
		32'h0000E108: begin
				q			<=			16'h3333;
		end
		32'h0000E10A: begin
				q			<=			16'h00B8;
		end
		32'h0000E10C: begin
				q			<=			16'h85B3;
		end
		32'h0000E10E: begin
				q			<=			16'h40E5;
		end
		32'h0000E110: begin
				q			<=			16'h2C23;
		end
		32'h0000E112: begin
				q			<=			16'h02B1;
		end
		32'h0000E114: begin
				q			<=			16'h0663;
		end
		32'h0000E116: begin
				q			<=			16'h0007;
		end
		32'h0000E118: begin
				q			<=			16'h88B3;
		end
		32'h0000E11A: begin
				q			<=			16'h4108;
		end
		32'h0000E11C: begin
				q			<=			16'hB693;
		end
		32'h0000E11E: begin
				q			<=			16'h0018;
		end
		32'h0000E120: begin
				q			<=			16'h2783;
		end
		32'h0000E122: begin
				q			<=			16'h02C1;
		end
		32'h0000E124: begin
				q			<=			16'hE8B3;
		end
		32'h0000E126: begin
				q			<=			16'h0066;
		end
		32'h0000E128: begin
				q			<=			16'h87B3;
		end
		32'h0000E12A: begin
				q			<=			16'h41D7;
		end
		32'h0000E12C: begin
				q			<=			16'h87B3;
		end
		32'h0000E12E: begin
				q			<=			16'h4117;
		end
		32'h0000E130: begin
				q			<=			16'h2E23;
		end
		32'h0000E132: begin
				q			<=			16'h02F1;
		end
		32'h0000E134: begin
				q			<=			16'h0413;
		end
		32'h0000E136: begin
				q			<=			16'h0006;
		end
		32'h0000E138: begin
				q			<=			16'h0913;
		end
		32'h0000E13A: begin
				q			<=			16'h0005;
		end
		32'h0000E13C: begin
				q			<=			16'hF06F;
		end
		32'h0000E13E: begin
				q			<=			16'hD49F;
		end
		32'h0000E140: begin
				q			<=			16'h86B7;
		end
		32'h0000E142: begin
				q			<=			16'h0000;
		end
		32'h0000E144: begin
				q			<=			16'h8693;
		end
		32'h0000E146: begin
				q			<=			16'hFFF6;
		end
		32'h0000E148: begin
				q			<=			16'h08E3;
		end
		32'h0000E14A: begin
				q			<=			16'hF4D6;
		end
		32'h0000E14C: begin
				q			<=			16'h4713;
		end
		32'h0000E14E: begin
				q			<=			16'hFFF7;
		end
		32'h0000E150: begin
				q			<=			16'h0793;
		end
		32'h0000E152: begin
				q			<=			16'h0740;
		end
		32'h0000E154: begin
				q			<=			16'hD263;
		end
		32'h0000E156: begin
				q			<=			16'h04E7;
		end
		32'h0000E158: begin
				q			<=			16'h0793;
		end
		32'h0000E15A: begin
				q			<=			16'h0010;
		end
		32'h0000E15C: begin
				q			<=			16'h2E23;
		end
		32'h0000E15E: begin
				q			<=			16'h0001;
		end
		32'h0000E160: begin
				q			<=			16'h2C23;
		end
		32'h0000E162: begin
				q			<=			16'h0001;
		end
		32'h0000E164: begin
				q			<=			16'h2A23;
		end
		32'h0000E166: begin
				q			<=			16'h0001;
		end
		32'h0000E168: begin
				q			<=			16'h2823;
		end
		32'h0000E16A: begin
				q			<=			16'h00F1;
		end
		32'h0000E16C: begin
				q			<=			16'h006F;
		end
		32'h0000E16E: begin
				q			<=			16'h0740;
		end
		32'h0000E170: begin
				q			<=			16'h86B7;
		end
		32'h0000E172: begin
				q			<=			16'h0000;
		end
		32'h0000E174: begin
				q			<=			16'h8693;
		end
		32'h0000E176: begin
				q			<=			16'hFFF6;
		end
		32'h0000E178: begin
				q			<=			16'h00E3;
		end
		32'h0000E17A: begin
				q			<=			16'hF2D6;
		end
		32'h0000E17C: begin
				q			<=			16'h2783;
		end
		32'h0000E17E: begin
				q			<=			16'h01C1;
		end
		32'h0000E180: begin
				q			<=			16'h06B7;
		end
		32'h0000E182: begin
				q			<=			16'h0008;
		end
		32'h0000E184: begin
				q			<=			16'hE7B3;
		end
		32'h0000E186: begin
				q			<=			16'h00D7;
		end
		32'h0000E188: begin
				q			<=			16'h2E23;
		end
		32'h0000E18A: begin
				q			<=			16'h00F1;
		end
		32'h0000E18C: begin
				q			<=			16'h0793;
		end
		32'h0000E18E: begin
				q			<=			16'hF8C0;
		end
		32'h0000E190: begin
				q			<=			16'h44E3;
		end
		32'h0000E192: begin
				q			<=			16'hFCF7;
		end
		32'h0000E194: begin
				q			<=			16'h0733;
		end
		32'h0000E196: begin
				q			<=			16'h40E0;
		end
		32'h0000E198: begin
				q			<=			16'h5693;
		end
		32'h0000E19A: begin
				q			<=			16'h4057;
		end
		32'h0000E19C: begin
				q			<=			16'h0893;
		end
		32'h0000E19E: begin
				q			<=			16'h0000;
		end
		32'h0000E1A0: begin
				q			<=			16'h7713;
		end
		32'h0000E1A2: begin
				q			<=			16'h01F7;
		end
		32'h0000E1A4: begin
				q			<=			16'h0793;
		end
		32'h0000E1A6: begin
				q			<=			16'h0000;
		end
		32'h0000E1A8: begin
				q			<=			16'h9313;
		end
		32'h0000E1AA: begin
				q			<=			16'h0027;
		end
		32'h0000E1AC: begin
				q			<=			16'h9663;
		end
		32'h0000E1AE: begin
				q			<=			16'h0AD7;
		end
		32'h0000E1B0: begin
				q			<=			16'h1A63;
		end
		32'h0000E1B2: begin
				q			<=			16'h0C07;
		end
		32'h0000E1B4: begin
				q			<=			16'h0693;
		end
		32'h0000E1B6: begin
				q			<=			16'h0030;
		end
		32'h0000E1B8: begin
				q			<=			16'h86B3;
		end
		32'h0000E1BA: begin
				q			<=			16'h40F6;
		end
		32'h0000E1BC: begin
				q			<=			16'hD863;
		end
		32'h0000E1BE: begin
				q			<=			16'h0AE6;
		end
		32'h0000E1C0: begin
				q			<=			16'h0713;
		end
		32'h0000E1C2: begin
				q			<=			16'h0040;
		end
		32'h0000E1C4: begin
				q			<=			16'h07B3;
		end
		32'h0000E1C6: begin
				q			<=			16'h40F7;
		end
		32'h0000E1C8: begin
				q			<=			16'h0693;
		end
		32'h0000E1CA: begin
				q			<=			16'h0040;
		end
		32'h0000E1CC: begin
				q			<=			16'h9863;
		end
		32'h0000E1CE: begin
				q			<=			16'h12D7;
		end
		32'h0000E1D0: begin
				q			<=			16'h2783;
		end
		32'h0000E1D2: begin
				q			<=			16'h0101;
		end
		32'h0000E1D4: begin
				q			<=			16'h38B3;
		end
		32'h0000E1D6: begin
				q			<=			16'h0110;
		end
		32'h0000E1D8: begin
				q			<=			16'hE8B3;
		end
		32'h0000E1DA: begin
				q			<=			16'h0117;
		end
		32'h0000E1DC: begin
				q			<=			16'h2823;
		end
		32'h0000E1DE: begin
				q			<=			16'h0111;
		end
		32'h0000E1E0: begin
				q			<=			16'h2683;
		end
		32'h0000E1E2: begin
				q			<=			16'h0241;
		end
		32'h0000E1E4: begin
				q			<=			16'h2803;
		end
		32'h0000E1E6: begin
				q			<=			16'h0201;
		end
		32'h0000E1E8: begin
				q			<=			16'h2703;
		end
		32'h0000E1EA: begin
				q			<=			16'h0101;
		end
		32'h0000E1EC: begin
				q			<=			16'h2783;
		end
		32'h0000E1EE: begin
				q			<=			16'h0141;
		end
		32'h0000E1F0: begin
				q			<=			16'h0733;
		end
		32'h0000E1F2: begin
				q			<=			16'h40E8;
		end
		32'h0000E1F4: begin
				q			<=			16'h87B3;
		end
		32'h0000E1F6: begin
				q			<=			16'h40F6;
		end
		32'h0000E1F8: begin
				q			<=			16'hB5B3;
		end
		32'h0000E1FA: begin
				q			<=			16'h00F6;
		end
		32'h0000E1FC: begin
				q			<=			16'h36B3;
		end
		32'h0000E1FE: begin
				q			<=			16'h00E8;
		end
		32'h0000E200: begin
				q			<=			16'h86B3;
		end
		32'h0000E202: begin
				q			<=			16'h40D7;
		end
		32'h0000E204: begin
				q			<=			16'h2A23;
		end
		32'h0000E206: begin
				q			<=			16'h02D1;
		end
		32'h0000E208: begin
				q			<=			16'h2823;
		end
		32'h0000E20A: begin
				q			<=			16'h02E1;
		end
		32'h0000E20C: begin
				q			<=			16'h0693;
		end
		32'h0000E20E: begin
				q			<=			16'h0000;
		end
		32'h0000E210: begin
				q			<=			16'h7463;
		end
		32'h0000E212: begin
				q			<=			16'h00E8;
		end
		32'h0000E214: begin
				q			<=			16'hB693;
		end
		32'h0000E216: begin
				q			<=			16'h0017;
		end
		32'h0000E218: begin
				q			<=			16'hE6B3;
		end
		32'h0000E21A: begin
				q			<=			16'h00B6;
		end
		32'h0000E21C: begin
				q			<=			16'h2703;
		end
		32'h0000E21E: begin
				q			<=			16'h0181;
		end
		32'h0000E220: begin
				q			<=			16'h2583;
		end
		32'h0000E222: begin
				q			<=			16'h0281;
		end
		32'h0000E224: begin
				q			<=			16'h8733;
		end
		32'h0000E226: begin
				q			<=			16'h40E5;
		end
		32'h0000E228: begin
				q			<=			16'h07B3;
		end
		32'h0000E22A: begin
				q			<=			16'h40D7;
		end
		32'h0000E22C: begin
				q			<=			16'h2C23;
		end
		32'h0000E22E: begin
				q			<=			16'h02F1;
		end
		32'h0000E230: begin
				q			<=			16'hB833;
		end
		32'h0000E232: begin
				q			<=			16'h00E5;
		end
		32'h0000E234: begin
				q			<=			16'h0593;
		end
		32'h0000E236: begin
				q			<=			16'h0000;
		end
		32'h0000E238: begin
				q			<=			16'h8463;
		end
		32'h0000E23A: begin
				q			<=			16'h0006;
		end
		32'h0000E23C: begin
				q			<=			16'h3593;
		end
		32'h0000E23E: begin
				q			<=			16'h0017;
		end
		32'h0000E240: begin
				q			<=			16'h2783;
		end
		32'h0000E242: begin
				q			<=			16'h02C1;
		end
		32'h0000E244: begin
				q			<=			16'h2703;
		end
		32'h0000E246: begin
				q			<=			16'h01C1;
		end
		32'h0000E248: begin
				q			<=			16'hE5B3;
		end
		32'h0000E24A: begin
				q			<=			16'h0105;
		end
		32'h0000E24C: begin
				q			<=			16'h87B3;
		end
		32'h0000E24E: begin
				q			<=			16'h40E7;
		end
		32'h0000E250: begin
				q			<=			16'h87B3;
		end
		32'h0000E252: begin
				q			<=			16'h40B7;
		end
		32'h0000E254: begin
				q			<=			16'hF06F;
		end
		32'h0000E256: begin
				q			<=			16'hEDDF;
		end
		32'h0000E258: begin
				q			<=			16'h0333;
		end
		32'h0000E25A: begin
				q			<=			16'h0068;
		end
		32'h0000E25C: begin
				q			<=			16'h2303;
		end
		32'h0000E25E: begin
				q			<=			16'h0003;
		end
		32'h0000E260: begin
				q			<=			16'h8793;
		end
		32'h0000E262: begin
				q			<=			16'h0017;
		end
		32'h0000E264: begin
				q			<=			16'hE8B3;
		end
		32'h0000E266: begin
				q			<=			16'h0068;
		end
		32'h0000E268: begin
				q			<=			16'hF06F;
		end
		32'h0000E26A: begin
				q			<=			16'hF41F;
		end
		32'h0000E26C: begin
				q			<=			16'h8E33;
		end
		32'h0000E26E: begin
				q			<=			16'h0065;
		end
		32'h0000E270: begin
				q			<=			16'h2E03;
		end
		32'h0000E272: begin
				q			<=			16'h000E;
		end
		32'h0000E274: begin
				q			<=			16'h0713;
		end
		32'h0000E276: begin
				q			<=			16'h0017;
		end
		32'h0000E278: begin
				q			<=			16'h8593;
		end
		32'h0000E27A: begin
				q			<=			16'h0045;
		end
		32'h0000E27C: begin
				q			<=			16'hAE23;
		end
		32'h0000E27E: begin
				q			<=			16'hFFC5;
		end
		32'h0000E280: begin
				q			<=			16'hF06F;
		end
		32'h0000E282: begin
				q			<=			16'hF3DF;
		end
		32'h0000E284: begin
				q			<=			16'h0693;
		end
		32'h0000E286: begin
				q			<=			16'h0401;
		end
		32'h0000E288: begin
				q			<=			16'h86B3;
		end
		32'h0000E28A: begin
				q			<=			16'h0066;
		end
		32'h0000E28C: begin
				q			<=			16'hA683;
		end
		32'h0000E28E: begin
				q			<=			16'hFD06;
		end
		32'h0000E290: begin
				q			<=			16'h0E93;
		end
		32'h0000E292: begin
				q			<=			16'h0200;
		end
		32'h0000E294: begin
				q			<=			16'h8EB3;
		end
		32'h0000E296: begin
				q			<=			16'h40EE;
		end
		32'h0000E298: begin
				q			<=			16'h96B3;
		end
		32'h0000E29A: begin
				q			<=			16'h01D6;
		end
		32'h0000E29C: begin
				q			<=			16'hE8B3;
		end
		32'h0000E29E: begin
				q			<=			16'h00D8;
		end
		32'h0000E2A0: begin
				q			<=			16'h0693;
		end
		32'h0000E2A2: begin
				q			<=			16'h0030;
		end
		32'h0000E2A4: begin
				q			<=			16'h0F13;
		end
		32'h0000E2A6: begin
				q			<=			16'h0000;
		end
		32'h0000E2A8: begin
				q			<=			16'h86B3;
		end
		32'h0000E2AA: begin
				q			<=			16'h40F6;
		end
		32'h0000E2AC: begin
				q			<=			16'h4463;
		end
		32'h0000E2AE: begin
				q			<=			16'h02DF;
		end
		32'h0000E2B0: begin
				q			<=			16'h0593;
		end
		32'h0000E2B2: begin
				q			<=			16'h0040;
		end
		32'h0000E2B4: begin
				q			<=			16'h87B3;
		end
		32'h0000E2B6: begin
				q			<=			16'h40F5;
		end
		32'h0000E2B8: begin
				q			<=			16'h9693;
		end
		32'h0000E2BA: begin
				q			<=			16'h0026;
		end
		32'h0000E2BC: begin
				q			<=			16'h0593;
		end
		32'h0000E2BE: begin
				q			<=			16'h0401;
		end
		32'h0000E2C0: begin
				q			<=			16'h86B3;
		end
		32'h0000E2C2: begin
				q			<=			16'h00D5;
		end
		32'h0000E2C4: begin
				q			<=			16'h2583;
		end
		32'h0000E2C6: begin
				q			<=			16'h01C1;
		end
		32'h0000E2C8: begin
				q			<=			16'hD733;
		end
		32'h0000E2CA: begin
				q			<=			16'h00E5;
		end
		32'h0000E2CC: begin
				q			<=			16'hA823;
		end
		32'h0000E2CE: begin
				q			<=			16'hFCE6;
		end
		32'h0000E2D0: begin
				q			<=			16'hF06F;
		end
		32'h0000E2D2: begin
				q			<=			16'hEF9F;
		end
		32'h0000E2D4: begin
				q			<=			16'h8FB3;
		end
		32'h0000E2D6: begin
				q			<=			16'h0065;
		end
		32'h0000E2D8: begin
				q			<=			16'hAE03;
		end
		32'h0000E2DA: begin
				q			<=			16'h000F;
		end
		32'h0000E2DC: begin
				q			<=			16'hAF83;
		end
		32'h0000E2DE: begin
				q			<=			16'h004F;
		end
		32'h0000E2E0: begin
				q			<=			16'h0F13;
		end
		32'h0000E2E2: begin
				q			<=			16'h001F;
		end
		32'h0000E2E4: begin
				q			<=			16'h5E33;
		end
		32'h0000E2E6: begin
				q			<=			16'h00EE;
		end
		32'h0000E2E8: begin
				q			<=			16'h9FB3;
		end
		32'h0000E2EA: begin
				q			<=			16'h01DF;
		end
		32'h0000E2EC: begin
				q			<=			16'h6E33;
		end
		32'h0000E2EE: begin
				q			<=			16'h01FE;
		end
		32'h0000E2F0: begin
				q			<=			16'hA023;
		end
		32'h0000E2F2: begin
				q			<=			16'h01C5;
		end
		32'h0000E2F4: begin
				q			<=			16'h8593;
		end
		32'h0000E2F6: begin
				q			<=			16'h0045;
		end
		32'h0000E2F8: begin
				q			<=			16'hF06F;
		end
		32'h0000E2FA: begin
				q			<=			16'hFB5F;
		end
		32'h0000E2FC: begin
				q			<=			16'h9713;
		end
		32'h0000E2FE: begin
				q			<=			16'h0027;
		end
		32'h0000E300: begin
				q			<=			16'h0733;
		end
		32'h0000E302: begin
				q			<=			16'h00E8;
		end
		32'h0000E304: begin
				q			<=			16'h2023;
		end
		32'h0000E306: begin
				q			<=			16'h0007;
		end
		32'h0000E308: begin
				q			<=			16'h8793;
		end
		32'h0000E30A: begin
				q			<=			16'h0017;
		end
		32'h0000E30C: begin
				q			<=			16'hF06F;
		end
		32'h0000E30E: begin
				q			<=			16'hEC1F;
		end
		32'h0000E310: begin
				q			<=			16'h8FB7;
		end
		32'h0000E312: begin
				q			<=			16'h0000;
		end
		32'h0000E314: begin
				q			<=			16'h0813;
		end
		32'h0000E316: begin
				q			<=			16'h0014;
		end
		32'h0000E318: begin
				q			<=			16'h8293;
		end
		32'h0000E31A: begin
				q			<=			16'hFFFF;
		end
		32'h0000E31C: begin
				q			<=			16'h7833;
		end
		32'h0000E31E: begin
				q			<=			16'h0058;
		end
		32'h0000E320: begin
				q			<=			16'h0F13;
		end
		32'h0000E322: begin
				q			<=			16'h0010;
		end
		32'h0000E324: begin
				q			<=			16'h2583;
		end
		32'h0000E326: begin
				q			<=			16'h0241;
		end
		32'h0000E328: begin
				q			<=			16'h2603;
		end
		32'h0000E32A: begin
				q			<=			16'h0141;
		end
		32'h0000E32C: begin
				q			<=			16'h2883;
		end
		32'h0000E32E: begin
				q			<=			16'h0181;
		end
		32'h0000E330: begin
				q			<=			16'h2E83;
		end
		32'h0000E332: begin
				q			<=			16'h01C1;
		end
		32'h0000E334: begin
				q			<=			16'h2303;
		end
		32'h0000E336: begin
				q			<=			16'h0281;
		end
		32'h0000E338: begin
				q			<=			16'h2E03;
		end
		32'h0000E33A: begin
				q			<=			16'h02C1;
		end
		32'h0000E33C: begin
				q			<=			16'h4E63;
		end
		32'h0000E33E: begin
				q			<=			16'h1D0F;
		end
		32'h0000E340: begin
				q			<=			16'hE833;
		end
		32'h0000E342: begin
				q			<=			16'h0065;
		end
		32'h0000E344: begin
				q			<=			16'h6F33;
		end
		32'h0000E346: begin
				q			<=			16'h0116;
		end
		32'h0000E348: begin
				q			<=			16'h6833;
		end
		32'h0000E34A: begin
				q			<=			16'h01C8;
		end
		32'h0000E34C: begin
				q			<=			16'h6F33;
		end
		32'h0000E34E: begin
				q			<=			16'h01DF;
		end
		32'h0000E350: begin
				q			<=			16'h6833;
		end
		32'h0000E352: begin
				q			<=			16'h00F8;
		end
		32'h0000E354: begin
				q			<=			16'h6F33;
		end
		32'h0000E356: begin
				q			<=			16'h00DF;
		end
		32'h0000E358: begin
				q			<=			16'h1863;
		end
		32'h0000E35A: begin
				q			<=			16'h1004;
		end
		32'h0000E35C: begin
				q			<=			16'h1263;
		end
		32'h0000E35E: begin
				q			<=			16'h020F;
		end
		32'h0000E360: begin
				q			<=			16'h2823;
		end
		32'h0000E362: begin
				q			<=			16'h02F1;
		end
		32'h0000E364: begin
				q			<=			16'h2A23;
		end
		32'h0000E366: begin
				q			<=			16'h02B1;
		end
		32'h0000E368: begin
				q			<=			16'h2C23;
		end
		32'h0000E36A: begin
				q			<=			16'h0261;
		end
		32'h0000E36C: begin
				q			<=			16'h2E23;
		end
		32'h0000E36E: begin
				q			<=			16'h03C1;
		end
		32'h0000E370: begin
				q			<=			16'h14E3;
		end
		32'h0000E372: begin
				q			<=			16'hD408;
		end
		32'h0000E374: begin
				q			<=			16'h0413;
		end
		32'h0000E376: begin
				q			<=			16'h0000;
		end
		32'h0000E378: begin
				q			<=			16'h0913;
		end
		32'h0000E37A: begin
				q			<=			16'h0000;
		end
		32'h0000E37C: begin
				q			<=			16'hF06F;
		end
		32'h0000E37E: begin
				q			<=			16'hD00F;
		end
		32'h0000E380: begin
				q			<=			16'h1C63;
		end
		32'h0000E382: begin
				q			<=			16'h0008;
		end
		32'h0000E384: begin
				q			<=			16'h2823;
		end
		32'h0000E386: begin
				q			<=			16'h02D1;
		end
		32'h0000E388: begin
				q			<=			16'h2A23;
		end
		32'h0000E38A: begin
				q			<=			16'h02C1;
		end
		32'h0000E38C: begin
				q			<=			16'h2C23;
		end
		32'h0000E38E: begin
				q			<=			16'h0311;
		end
		32'h0000E390: begin
				q			<=			16'h2E23;
		end
		32'h0000E392: begin
				q			<=			16'h03D1;
		end
		32'h0000E394: begin
				q			<=			16'hF06F;
		end
		32'h0000E396: begin
				q			<=			16'hC98F;
		end
		32'h0000E398: begin
				q			<=			16'h8833;
		end
		32'h0000E39A: begin
				q			<=			16'h40F6;
		end
		32'h0000E39C: begin
				q			<=			16'h02B3;
		end
		32'h0000E39E: begin
				q			<=			16'h40B6;
		end
		32'h0000E3A0: begin
				q			<=			16'hBFB3;
		end
		32'h0000E3A2: begin
				q			<=			16'h0106;
		end
		32'h0000E3A4: begin
				q			<=			16'h3F33;
		end
		32'h0000E3A6: begin
				q			<=			16'h0056;
		end
		32'h0000E3A8: begin
				q			<=			16'h82B3;
		end
		32'h0000E3AA: begin
				q			<=			16'h41F2;
		end
		32'h0000E3AC: begin
				q			<=			16'h2823;
		end
		32'h0000E3AE: begin
				q			<=			16'h0301;
		end
		32'h0000E3B0: begin
				q			<=			16'h2A23;
		end
		32'h0000E3B2: begin
				q			<=			16'h0251;
		end
		32'h0000E3B4: begin
				q			<=			16'h0F93;
		end
		32'h0000E3B6: begin
				q			<=			16'h0000;
		end
		32'h0000E3B8: begin
				q			<=			16'hF663;
		end
		32'h0000E3BA: begin
				q			<=			16'h0106;
		end
		32'h0000E3BC: begin
				q			<=			16'h8FB3;
		end
		32'h0000E3BE: begin
				q			<=			16'h40C5;
		end
		32'h0000E3C0: begin
				q			<=			16'hBF93;
		end
		32'h0000E3C2: begin
				q			<=			16'h001F;
		end
		32'h0000E3C4: begin
				q			<=			16'h83B3;
		end
		32'h0000E3C6: begin
				q			<=			16'h4068;
		end
		32'h0000E3C8: begin
				q			<=			16'hEFB3;
		end
		32'h0000E3CA: begin
				q			<=			16'h01EF;
		end
		32'h0000E3CC: begin
				q			<=			16'h8A33;
		end
		32'h0000E3CE: begin
				q			<=			16'h41F3;
		end
		32'h0000E3D0: begin
				q			<=			16'h2C23;
		end
		32'h0000E3D2: begin
				q			<=			16'h0341;
		end
		32'h0000E3D4: begin
				q			<=			16'hBAB3;
		end
		32'h0000E3D6: begin
				q			<=			16'h0078;
		end
		32'h0000E3D8: begin
				q			<=			16'h0993;
		end
		32'h0000E3DA: begin
				q			<=			16'h0000;
		end
		32'h0000E3DC: begin
				q			<=			16'h8463;
		end
		32'h0000E3DE: begin
				q			<=			16'h000F;
		end
		32'h0000E3E0: begin
				q			<=			16'hB993;
		end
		32'h0000E3E2: begin
				q			<=			16'h0013;
		end
		32'h0000E3E4: begin
				q			<=			16'h8F33;
		end
		32'h0000E3E6: begin
				q			<=			16'h41CE;
		end
		32'h0000E3E8: begin
				q			<=			16'hE9B3;
		end
		32'h0000E3EA: begin
				q			<=			16'h0159;
		end
		32'h0000E3EC: begin
				q			<=			16'h0F33;
		end
		32'h0000E3EE: begin
				q			<=			16'h413F;
		end
		32'h0000E3F0: begin
				q			<=			16'h2E23;
		end
		32'h0000E3F2: begin
				q			<=			16'h03E1;
		end
		32'h0000E3F4: begin
				q			<=			16'h1F93;
		end
		32'h0000E3F6: begin
				q			<=			16'h00CF;
		end
		32'h0000E3F8: begin
				q			<=			16'hDE63;
		end
		32'h0000E3FA: begin
				q			<=			16'h040F;
		end
		32'h0000E3FC: begin
				q			<=			16'h86B3;
		end
		32'h0000E3FE: begin
				q			<=			16'h40D7;
		end
		32'h0000E400: begin
				q			<=			16'h8633;
		end
		32'h0000E402: begin
				q			<=			16'h40C5;
		end
		32'h0000E404: begin
				q			<=			16'hB833;
		end
		32'h0000E406: begin
				q			<=			16'h00D7;
		end
		32'h0000E408: begin
				q			<=			16'h0833;
		end
		32'h0000E40A: begin
				q			<=			16'h4106;
		end
		32'h0000E40C: begin
				q			<=			16'h2A23;
		end
		32'h0000E40E: begin
				q			<=			16'h0301;
		end
		32'h0000E410: begin
				q			<=			16'h2823;
		end
		32'h0000E412: begin
				q			<=			16'h02D1;
		end
		32'h0000E414: begin
				q			<=			16'hB5B3;
		end
		32'h0000E416: begin
				q			<=			16'h00C5;
		end
		32'h0000E418: begin
				q			<=			16'h0813;
		end
		32'h0000E41A: begin
				q			<=			16'h0000;
		end
		32'h0000E41C: begin
				q			<=			16'hF463;
		end
		32'h0000E41E: begin
				q			<=			16'h00D7;
		end
		32'h0000E420: begin
				q			<=			16'h3813;
		end
		32'h0000E422: begin
				q			<=			16'h0016;
		end
		32'h0000E424: begin
				q			<=			16'h07B3;
		end
		32'h0000E426: begin
				q			<=			16'h4113;
		end
		32'h0000E428: begin
				q			<=			16'h65B3;
		end
		32'h0000E42A: begin
				q			<=			16'h00B8;
		end
		32'h0000E42C: begin
				q			<=			16'h36B3;
		end
		32'h0000E42E: begin
				q			<=			16'h00F3;
		end
		32'h0000E430: begin
				q			<=			16'h87B3;
		end
		32'h0000E432: begin
				q			<=			16'h40B7;
		end
		32'h0000E434: begin
				q			<=			16'h2C23;
		end
		32'h0000E436: begin
				q			<=			16'h02F1;
		end
		32'h0000E438: begin
				q			<=			16'h8463;
		end
		32'h0000E43A: begin
				q			<=			16'h0005;
		end
		32'h0000E43C: begin
				q			<=			16'hB713;
		end
		32'h0000E43E: begin
				q			<=			16'h0013;
		end
		32'h0000E440: begin
				q			<=			16'h07B3;
		end
		32'h0000E442: begin
				q			<=			16'h41DE;
		end
		32'h0000E444: begin
				q			<=			16'h6733;
		end
		32'h0000E446: begin
				q			<=			16'h00D7;
		end
		32'h0000E448: begin
				q			<=			16'h8733;
		end
		32'h0000E44A: begin
				q			<=			16'h40E7;
		end
		32'h0000E44C: begin
				q			<=			16'h2E23;
		end
		32'h0000E44E: begin
				q			<=			16'h02E1;
		end
		32'h0000E450: begin
				q			<=			16'hF06F;
		end
		32'h0000E452: begin
				q			<=			16'hC69F;
		end
		32'h0000E454: begin
				q			<=			16'h6833;
		end
		32'h0000E456: begin
				q			<=			16'h0058;
		end
		32'h0000E458: begin
				q			<=			16'h6833;
		end
		32'h0000E45A: begin
				q			<=			16'h0148;
		end
		32'h0000E45C: begin
				q			<=			16'h6833;
		end
		32'h0000E45E: begin
				q			<=			16'h01E8;
		end
		32'h0000E460: begin
				q			<=			16'h0AE3;
		end
		32'h0000E462: begin
				q			<=			16'hF008;
		end
		32'h0000E464: begin
				q			<=			16'hF06F;
		end
		32'h0000E466: begin
				q			<=			16'hBC8F;
		end
		32'h0000E468: begin
				q			<=			16'h0393;
		end
		32'h0000E46A: begin
				q			<=			16'h0301;
		end
		32'h0000E46C: begin
				q			<=			16'h1E63;
		end
		32'h0000E46E: begin
				q			<=			16'h040F;
		end
		32'h0000E470: begin
				q			<=			16'h1E63;
		end
		32'h0000E472: begin
				q			<=			16'h0208;
		end
		32'h0000E474: begin
				q			<=			16'h2E23;
		end
		32'h0000E476: begin
				q			<=			16'h03F1;
		end
		32'h0000E478: begin
				q			<=			16'h2C23;
		end
		32'h0000E47A: begin
				q			<=			16'h0201;
		end
		32'h0000E47C: begin
				q			<=			16'h2A23;
		end
		32'h0000E47E: begin
				q			<=			16'h0201;
		end
		32'h0000E480: begin
				q			<=			16'h2823;
		end
		32'h0000E482: begin
				q			<=			16'h0201;
		end
		32'h0000E484: begin
				q			<=			16'h0793;
		end
		32'h0000E486: begin
				q			<=			16'h03C1;
		end
		32'h0000E488: begin
				q			<=			16'hA703;
		end
		32'h0000E48A: begin
				q			<=			16'h0007;
		end
		32'h0000E48C: begin
				q			<=			16'hA683;
		end
		32'h0000E48E: begin
				q			<=			16'hFFC7;
		end
		32'h0000E490: begin
				q			<=			16'h8793;
		end
		32'h0000E492: begin
				q			<=			16'hFFC7;
		end
		32'h0000E494: begin
				q			<=			16'h1713;
		end
		32'h0000E496: begin
				q			<=			16'h0037;
		end
		32'h0000E498: begin
				q			<=			16'hD693;
		end
		32'h0000E49A: begin
				q			<=			16'h01D6;
		end
		32'h0000E49C: begin
				q			<=			16'h6733;
		end
		32'h0000E49E: begin
				q			<=			16'h00D7;
		end
		32'h0000E4A0: begin
				q			<=			16'hA223;
		end
		32'h0000E4A2: begin
				q			<=			16'h00E7;
		end
		32'h0000E4A4: begin
				q			<=			16'h92E3;
		end
		32'h0000E4A6: begin
				q			<=			16'hFEF3;
		end
		32'h0000E4A8: begin
				q			<=			16'hF06F;
		end
		32'h0000E4AA: begin
				q			<=			16'h881F;
		end
		32'h0000E4AC: begin
				q			<=			16'h2823;
		end
		32'h0000E4AE: begin
				q			<=			16'h02F1;
		end
		32'h0000E4B0: begin
				q			<=			16'h2A23;
		end
		32'h0000E4B2: begin
				q			<=			16'h02B1;
		end
		32'h0000E4B4: begin
				q			<=			16'h2C23;
		end
		32'h0000E4B6: begin
				q			<=			16'h0261;
		end
		32'h0000E4B8: begin
				q			<=			16'h2E23;
		end
		32'h0000E4BA: begin
				q			<=			16'h03C1;
		end
		32'h0000E4BC: begin
				q			<=			16'h0913;
		end
		32'h0000E4BE: begin
				q			<=			16'h0005;
		end
		32'h0000E4C0: begin
				q			<=			16'h8413;
		end
		32'h0000E4C2: begin
				q			<=			16'h0002;
		end
		32'h0000E4C4: begin
				q			<=			16'hF06F;
		end
		32'h0000E4C6: begin
				q			<=			16'hB68F;
		end
		32'h0000E4C8: begin
				q			<=			16'h1C63;
		end
		32'h0000E4CA: begin
				q			<=			16'h0008;
		end
		32'h0000E4CC: begin
				q			<=			16'h2823;
		end
		32'h0000E4CE: begin
				q			<=			16'h02D1;
		end
		32'h0000E4D0: begin
				q			<=			16'h2A23;
		end
		32'h0000E4D2: begin
				q			<=			16'h02C1;
		end
		32'h0000E4D4: begin
				q			<=			16'h2C23;
		end
		32'h0000E4D6: begin
				q			<=			16'h0311;
		end
		32'h0000E4D8: begin
				q			<=			16'h2E23;
		end
		32'h0000E4DA: begin
				q			<=			16'h03D1;
		end
		32'h0000E4DC: begin
				q			<=			16'hF06F;
		end
		32'h0000E4DE: begin
				q			<=			16'hFE5F;
		end
		32'h0000E4E0: begin
				q			<=			16'h2E23;
		end
		32'h0000E4E2: begin
				q			<=			16'h03F1;
		end
		32'h0000E4E4: begin
				q			<=			16'h2C23;
		end
		32'h0000E4E6: begin
				q			<=			16'h0201;
		end
		32'h0000E4E8: begin
				q			<=			16'h2A23;
		end
		32'h0000E4EA: begin
				q			<=			16'h0201;
		end
		32'h0000E4EC: begin
				q			<=			16'h2823;
		end
		32'h0000E4EE: begin
				q			<=			16'h0201;
		end
		32'h0000E4F0: begin
				q			<=			16'h0793;
		end
		32'h0000E4F2: begin
				q			<=			16'h03C1;
		end
		32'h0000E4F4: begin
				q			<=			16'hA703;
		end
		32'h0000E4F6: begin
				q			<=			16'h0007;
		end
		32'h0000E4F8: begin
				q			<=			16'hA683;
		end
		32'h0000E4FA: begin
				q			<=			16'hFFC7;
		end
		32'h0000E4FC: begin
				q			<=			16'h8793;
		end
		32'h0000E4FE: begin
				q			<=			16'hFFC7;
		end
		32'h0000E500: begin
				q			<=			16'h1713;
		end
		32'h0000E502: begin
				q			<=			16'h0037;
		end
		32'h0000E504: begin
				q			<=			16'hD693;
		end
		32'h0000E506: begin
				q			<=			16'h01D6;
		end
		32'h0000E508: begin
				q			<=			16'h6733;
		end
		32'h0000E50A: begin
				q			<=			16'h00D7;
		end
		32'h0000E50C: begin
				q			<=			16'hA223;
		end
		32'h0000E50E: begin
				q			<=			16'h00E7;
		end
		32'h0000E510: begin
				q			<=			16'h92E3;
		end
		32'h0000E512: begin
				q			<=			16'hFEF3;
		end
		32'h0000E514: begin
				q			<=			16'hF06F;
		end
		32'h0000E516: begin
				q			<=			16'h815F;
		end
		32'h0000E518: begin
				q			<=			16'h8833;
		end
		32'h0000E51A: begin
				q			<=			16'h40F6;
		end
		32'h0000E51C: begin
				q			<=			16'h02B3;
		end
		32'h0000E51E: begin
				q			<=			16'h40B6;
		end
		32'h0000E520: begin
				q			<=			16'hBFB3;
		end
		32'h0000E522: begin
				q			<=			16'h0106;
		end
		32'h0000E524: begin
				q			<=			16'h3F33;
		end
		32'h0000E526: begin
				q			<=			16'h0056;
		end
		32'h0000E528: begin
				q			<=			16'h82B3;
		end
		32'h0000E52A: begin
				q			<=			16'h41F2;
		end
		32'h0000E52C: begin
				q			<=			16'h2823;
		end
		32'h0000E52E: begin
				q			<=			16'h0301;
		end
		32'h0000E530: begin
				q			<=			16'h2A23;
		end
		32'h0000E532: begin
				q			<=			16'h0251;
		end
		32'h0000E534: begin
				q			<=			16'h0F93;
		end
		32'h0000E536: begin
				q			<=			16'h0000;
		end
		32'h0000E538: begin
				q			<=			16'hF663;
		end
		32'h0000E53A: begin
				q			<=			16'h0106;
		end
		32'h0000E53C: begin
				q			<=			16'h8FB3;
		end
		32'h0000E53E: begin
				q			<=			16'h40C5;
		end
		32'h0000E540: begin
				q			<=			16'hBF93;
		end
		32'h0000E542: begin
				q			<=			16'h001F;
		end
		32'h0000E544: begin
				q			<=			16'h83B3;
		end
		32'h0000E546: begin
				q			<=			16'h4068;
		end
		32'h0000E548: begin
				q			<=			16'hEFB3;
		end
		32'h0000E54A: begin
				q			<=			16'h01EF;
		end
		32'h0000E54C: begin
				q			<=			16'h8A33;
		end
		32'h0000E54E: begin
				q			<=			16'h41F3;
		end
		32'h0000E550: begin
				q			<=			16'h2C23;
		end
		32'h0000E552: begin
				q			<=			16'h0341;
		end
		32'h0000E554: begin
				q			<=			16'hBAB3;
		end
		32'h0000E556: begin
				q			<=			16'h0078;
		end
		32'h0000E558: begin
				q			<=			16'h0993;
		end
		32'h0000E55A: begin
				q			<=			16'h0000;
		end
		32'h0000E55C: begin
				q			<=			16'h8463;
		end
		32'h0000E55E: begin
				q			<=			16'h000F;
		end
		32'h0000E560: begin
				q			<=			16'hB993;
		end
		32'h0000E562: begin
				q			<=			16'h0013;
		end
		32'h0000E564: begin
				q			<=			16'h8F33;
		end
		32'h0000E566: begin
				q			<=			16'h41CE;
		end
		32'h0000E568: begin
				q			<=			16'hE9B3;
		end
		32'h0000E56A: begin
				q			<=			16'h0159;
		end
		32'h0000E56C: begin
				q			<=			16'h0F33;
		end
		32'h0000E56E: begin
				q			<=			16'h413F;
		end
		32'h0000E570: begin
				q			<=			16'h2E23;
		end
		32'h0000E572: begin
				q			<=			16'h03E1;
		end
		32'h0000E574: begin
				q			<=			16'h1F93;
		end
		32'h0000E576: begin
				q			<=			16'h00CF;
		end
		32'h0000E578: begin
				q			<=			16'hDA63;
		end
		32'h0000E57A: begin
				q			<=			16'h0A0F;
		end
		32'h0000E57C: begin
				q			<=			16'h86B3;
		end
		32'h0000E57E: begin
				q			<=			16'h40D7;
		end
		32'h0000E580: begin
				q			<=			16'h8633;
		end
		32'h0000E582: begin
				q			<=			16'h40C5;
		end
		32'h0000E584: begin
				q			<=			16'hB833;
		end
		32'h0000E586: begin
				q			<=			16'h00D7;
		end
		32'h0000E588: begin
				q			<=			16'h0833;
		end
		32'h0000E58A: begin
				q			<=			16'h4106;
		end
		32'h0000E58C: begin
				q			<=			16'h2A23;
		end
		32'h0000E58E: begin
				q			<=			16'h0301;
		end
		32'h0000E590: begin
				q			<=			16'h2823;
		end
		32'h0000E592: begin
				q			<=			16'h02D1;
		end
		32'h0000E594: begin
				q			<=			16'hB5B3;
		end
		32'h0000E596: begin
				q			<=			16'h00C5;
		end
		32'h0000E598: begin
				q			<=			16'h0813;
		end
		32'h0000E59A: begin
				q			<=			16'h0000;
		end
		32'h0000E59C: begin
				q			<=			16'hF463;
		end
		32'h0000E59E: begin
				q			<=			16'h00D7;
		end
		32'h0000E5A0: begin
				q			<=			16'h3813;
		end
		32'h0000E5A2: begin
				q			<=			16'h0016;
		end
		32'h0000E5A4: begin
				q			<=			16'h07B3;
		end
		32'h0000E5A6: begin
				q			<=			16'h4113;
		end
		32'h0000E5A8: begin
				q			<=			16'h65B3;
		end
		32'h0000E5AA: begin
				q			<=			16'h00B8;
		end
		32'h0000E5AC: begin
				q			<=			16'h36B3;
		end
		32'h0000E5AE: begin
				q			<=			16'h00F3;
		end
		32'h0000E5B0: begin
				q			<=			16'h87B3;
		end
		32'h0000E5B2: begin
				q			<=			16'h40B7;
		end
		32'h0000E5B4: begin
				q			<=			16'h2C23;
		end
		32'h0000E5B6: begin
				q			<=			16'h02F1;
		end
		32'h0000E5B8: begin
				q			<=			16'h8463;
		end
		32'h0000E5BA: begin
				q			<=			16'h0005;
		end
		32'h0000E5BC: begin
				q			<=			16'hB713;
		end
		32'h0000E5BE: begin
				q			<=			16'h0013;
		end
		32'h0000E5C0: begin
				q			<=			16'h07B3;
		end
		32'h0000E5C2: begin
				q			<=			16'h41DE;
		end
		32'h0000E5C4: begin
				q			<=			16'h6733;
		end
		32'h0000E5C6: begin
				q			<=			16'h00D7;
		end
		32'h0000E5C8: begin
				q			<=			16'h8733;
		end
		32'h0000E5CA: begin
				q			<=			16'h40E7;
		end
		32'h0000E5CC: begin
				q			<=			16'h2E23;
		end
		32'h0000E5CE: begin
				q			<=			16'h02E1;
		end
		32'h0000E5D0: begin
				q			<=			16'h0913;
		end
		32'h0000E5D2: begin
				q			<=			16'h0005;
		end
		32'h0000E5D4: begin
				q			<=			16'h2503;
		end
		32'h0000E5D6: begin
				q			<=			16'h03C1;
		end
		32'h0000E5D8: begin
				q			<=			16'h0463;
		end
		32'h0000E5DA: begin
				q			<=			16'h0605;
		end
		32'h0000E5DC: begin
				q			<=			16'h00EF;
		end
		32'h0000E5DE: begin
				q			<=			16'h2F10;
		end
		32'h0000E5E0: begin
				q			<=			16'h0513;
		end
		32'h0000E5E2: begin
				q			<=			16'hFF45;
		end
		32'h0000E5E4: begin
				q			<=			16'h0693;
		end
		32'h0000E5E6: begin
				q			<=			16'h0200;
		end
		32'h0000E5E8: begin
				q			<=			16'h6833;
		end
		32'h0000E5EA: begin
				q			<=			16'h02D5;
		end
		32'h0000E5EC: begin
				q			<=			16'h47B3;
		end
		32'h0000E5EE: begin
				q			<=			16'h02D5;
		end
		32'h0000E5F0: begin
				q			<=			16'h0463;
		end
		32'h0000E5F2: begin
				q			<=			16'h0808;
		end
		32'h0000E5F4: begin
				q			<=			16'h0713;
		end
		32'h0000E5F6: begin
				q			<=			16'hFFC0;
		end
		32'h0000E5F8: begin
				q			<=			16'h9593;
		end
		32'h0000E5FA: begin
				q			<=			16'h0027;
		end
		32'h0000E5FC: begin
				q			<=			16'h0E13;
		end
		32'h0000E5FE: begin
				q			<=			16'hFF00;
		end
		32'h0000E600: begin
				q			<=			16'h86B3;
		end
		32'h0000E602: begin
				q			<=			16'h4106;
		end
		32'h0000E604: begin
				q			<=			16'h8733;
		end
		32'h0000E606: begin
				q			<=			16'h02E7;
		end
		32'h0000E608: begin
				q			<=			16'h0713;
		end
		32'h0000E60A: begin
				q			<=			16'hFFC7;
		end
		32'h0000E60C: begin
				q			<=			16'h1863;
		end
		32'h0000E60E: begin
				q			<=			16'h11C7;
		end
		32'h0000E610: begin
				q			<=			16'h0713;
		end
		32'h0000E612: begin
				q			<=			16'h0401;
		end
		32'h0000E614: begin
				q			<=			16'h05B3;
		end
		32'h0000E616: begin
				q			<=			16'h00B7;
		end
		32'h0000E618: begin
				q			<=			16'h2703;
		end
		32'h0000E61A: begin
				q			<=			16'h0301;
		end
		32'h0000E61C: begin
				q			<=			16'h8793;
		end
		32'h0000E61E: begin
				q			<=			16'hFFF7;
		end
		32'h0000E620: begin
				q			<=			16'h1833;
		end
		32'h0000E622: begin
				q			<=			16'h0107;
		end
		32'h0000E624: begin
				q			<=			16'hA823;
		end
		32'h0000E626: begin
				q			<=			16'hFF05;
		end
		32'h0000E628: begin
				q			<=			16'h006F;
		end
		32'h0000E62A: begin
				q			<=			16'h07C0;
		end
		32'h0000E62C: begin
				q			<=			16'h6833;
		end
		32'h0000E62E: begin
				q			<=			16'h0058;
		end
		32'h0000E630: begin
				q			<=			16'h6833;
		end
		32'h0000E632: begin
				q			<=			16'h0148;
		end
		32'h0000E634: begin
				q			<=			16'h6833;
		end
		32'h0000E636: begin
				q			<=			16'h01E8;
		end
		32'h0000E638: begin
				q			<=			16'h0EE3;
		end
		32'h0000E63A: begin
				q			<=			16'hD208;
		end
		32'h0000E63C: begin
				q			<=			16'hF06F;
		end
		32'h0000E63E: begin
				q			<=			16'hF99F;
		end
		32'h0000E640: begin
				q			<=			16'h2503;
		end
		32'h0000E642: begin
				q			<=			16'h0381;
		end
		32'h0000E644: begin
				q			<=			16'h0863;
		end
		32'h0000E646: begin
				q			<=			16'h0005;
		end
		32'h0000E648: begin
				q			<=			16'h00EF;
		end
		32'h0000E64A: begin
				q			<=			16'h2850;
		end
		32'h0000E64C: begin
				q			<=			16'h0513;
		end
		32'h0000E64E: begin
				q			<=			16'h0205;
		end
		32'h0000E650: begin
				q			<=			16'hF06F;
		end
		32'h0000E652: begin
				q			<=			16'hF91F;
		end
		32'h0000E654: begin
				q			<=			16'h2503;
		end
		32'h0000E656: begin
				q			<=			16'h0341;
		end
		32'h0000E658: begin
				q			<=			16'h0863;
		end
		32'h0000E65A: begin
				q			<=			16'h0005;
		end
		32'h0000E65C: begin
				q			<=			16'h00EF;
		end
		32'h0000E65E: begin
				q			<=			16'h2710;
		end
		32'h0000E660: begin
				q			<=			16'h0513;
		end
		32'h0000E662: begin
				q			<=			16'h0405;
		end
		32'h0000E664: begin
				q			<=			16'hF06F;
		end
		32'h0000E666: begin
				q			<=			16'hF7DF;
		end
		32'h0000E668: begin
				q			<=			16'h2503;
		end
		32'h0000E66A: begin
				q			<=			16'h0301;
		end
		32'h0000E66C: begin
				q			<=			16'h00EF;
		end
		32'h0000E66E: begin
				q			<=			16'h2610;
		end
		32'h0000E670: begin
				q			<=			16'h0513;
		end
		32'h0000E672: begin
				q			<=			16'h0605;
		end
		32'h0000E674: begin
				q			<=			16'hF06F;
		end
		32'h0000E676: begin
				q			<=			16'hF6DF;
		end
		32'h0000E678: begin
				q			<=			16'h0613;
		end
		32'h0000E67A: begin
				q			<=			16'hFFC0;
		end
		32'h0000E67C: begin
				q			<=			16'h8633;
		end
		32'h0000E67E: begin
				q			<=			16'h02C7;
		end
		32'h0000E680: begin
				q			<=			16'h0713;
		end
		32'h0000E682: begin
				q			<=			16'h0301;
		end
		32'h0000E684: begin
				q			<=			16'h0693;
		end
		32'h0000E686: begin
				q			<=			16'h0030;
		end
		32'h0000E688: begin
				q			<=			16'h05B3;
		end
		32'h0000E68A: begin
				q			<=			16'h00C7;
		end
		32'h0000E68C: begin
				q			<=			16'hA583;
		end
		32'h0000E68E: begin
				q			<=			16'h00C5;
		end
		32'h0000E690: begin
				q			<=			16'h8693;
		end
		32'h0000E692: begin
				q			<=			16'hFFF6;
		end
		32'h0000E694: begin
				q			<=			16'h0713;
		end
		32'h0000E696: begin
				q			<=			16'hFFC7;
		end
		32'h0000E698: begin
				q			<=			16'h2823;
		end
		32'h0000E69A: begin
				q			<=			16'h00B7;
		end
		32'h0000E69C: begin
				q			<=			16'hD6E3;
		end
		32'h0000E69E: begin
				q			<=			16'hFEF6;
		end
		32'h0000E6A0: begin
				q			<=			16'h8793;
		end
		32'h0000E6A2: begin
				q			<=			16'hFFF7;
		end
		32'h0000E6A4: begin
				q			<=			16'h0693;
		end
		32'h0000E6A6: begin
				q			<=			16'hFFF0;
		end
		32'h0000E6A8: begin
				q			<=			16'h9063;
		end
		32'h0000E6AA: begin
				q			<=			16'h0AD7;
		end
		32'h0000E6AC: begin
				q			<=			16'h4063;
		end
		32'h0000E6AE: begin
				q			<=			16'h1885;
		end
		32'h0000E6B0: begin
				q			<=			16'h0433;
		end
		32'h0000E6B2: begin
				q			<=			16'h4085;
		end
		32'h0000E6B4: begin
				q			<=			16'h0713;
		end
		32'h0000E6B6: begin
				q			<=			16'h0200;
		end
		32'h0000E6B8: begin
				q			<=			16'h0413;
		end
		32'h0000E6BA: begin
				q			<=			16'h0014;
		end
		32'h0000E6BC: begin
				q			<=			16'h47B3;
		end
		32'h0000E6BE: begin
				q			<=			16'h02E4;
		end
		32'h0000E6C0: begin
				q			<=			16'h0513;
		end
		32'h0000E6C2: begin
				q			<=			16'h0000;
		end
		32'h0000E6C4: begin
				q			<=			16'h6433;
		end
		32'h0000E6C6: begin
				q			<=			16'h02E4;
		end
		32'h0000E6C8: begin
				q			<=			16'h0713;
		end
		32'h0000E6CA: begin
				q			<=			16'h0000;
		end
		32'h0000E6CC: begin
				q			<=			16'h4A63;
		end
		32'h0000E6CE: begin
				q			<=			16'h08F7;
		end
		32'h0000E6D0: begin
				q			<=			16'h8713;
		end
		32'h0000E6D2: begin
				q			<=			16'h0007;
		end
		32'h0000E6D4: begin
				q			<=			16'hD463;
		end
		32'h0000E6D6: begin
				q			<=			16'h0007;
		end
		32'h0000E6D8: begin
				q			<=			16'h0713;
		end
		32'h0000E6DA: begin
				q			<=			16'h0000;
		end
		32'h0000E6DC: begin
				q			<=			16'h9313;
		end
		32'h0000E6DE: begin
				q			<=			16'h0027;
		end
		32'h0000E6E0: begin
				q			<=			16'h1A63;
		end
		32'h0000E6E2: begin
				q			<=			16'h0A04;
		end
		32'h0000E6E4: begin
				q			<=			16'h0693;
		end
		32'h0000E6E6: begin
				q			<=			16'h0030;
		end
		32'h0000E6E8: begin
				q			<=			16'h0713;
		end
		32'h0000E6EA: begin
				q			<=			16'h0301;
		end
		32'h0000E6EC: begin
				q			<=			16'h86B3;
		end
		32'h0000E6EE: begin
				q			<=			16'h40F6;
		end
		32'h0000E6F0: begin
				q			<=			16'hD663;
		end
		32'h0000E6F2: begin
				q			<=			16'h0886;
		end
		32'h0000E6F4: begin
				q			<=			16'h0713;
		end
		32'h0000E6F6: begin
				q			<=			16'h0040;
		end
		32'h0000E6F8: begin
				q			<=			16'h07B3;
		end
		32'h0000E6FA: begin
				q			<=			16'h40F7;
		end
		32'h0000E6FC: begin
				q			<=			16'h0693;
		end
		32'h0000E6FE: begin
				q			<=			16'h0030;
		end
		32'h0000E700: begin
				q			<=			16'hDA63;
		end
		32'h0000E702: begin
				q			<=			16'h10F6;
		end
		32'h0000E704: begin
				q			<=			16'h2703;
		end
		32'h0000E706: begin
				q			<=			16'h0301;
		end
		32'h0000E708: begin
				q			<=			16'h37B3;
		end
		32'h0000E70A: begin
				q			<=			16'h00A0;
		end
		32'h0000E70C: begin
				q			<=			16'h0413;
		end
		32'h0000E70E: begin
				q			<=			16'h0000;
		end
		32'h0000E710: begin
				q			<=			16'h67B3;
		end
		32'h0000E712: begin
				q			<=			16'h00F7;
		end
		32'h0000E714: begin
				q			<=			16'h2823;
		end
		32'h0000E716: begin
				q			<=			16'h02F1;
		end
		32'h0000E718: begin
				q			<=			16'hF06F;
		end
		32'h0000E71A: begin
				q			<=			16'h914F;
		end
		32'h0000E71C: begin
				q			<=			16'h0613;
		end
		32'h0000E71E: begin
				q			<=			16'h0301;
		end
		32'h0000E720: begin
				q			<=			16'h0333;
		end
		32'h0000E722: begin
				q			<=			16'h00E6;
		end
		32'h0000E724: begin
				q			<=			16'h88B3;
		end
		32'h0000E726: begin
				q			<=			16'h00E5;
		end
		32'h0000E728: begin
				q			<=			16'h08B3;
		end
		32'h0000E72A: begin
				q			<=			16'h0116;
		end
		32'h0000E72C: begin
				q			<=			16'h2603;
		end
		32'h0000E72E: begin
				q			<=			16'h00C3;
		end
		32'h0000E730: begin
				q			<=			16'h2303;
		end
		32'h0000E732: begin
				q			<=			16'h0103;
		end
		32'h0000E734: begin
				q			<=			16'h5633;
		end
		32'h0000E736: begin
				q			<=			16'h00D6;
		end
		32'h0000E738: begin
				q			<=			16'h1333;
		end
		32'h0000E73A: begin
				q			<=			16'h0103;
		end
		32'h0000E73C: begin
				q			<=			16'h6633;
		end
		32'h0000E73E: begin
				q			<=			16'h0066;
		end
		32'h0000E740: begin
				q			<=			16'hA823;
		end
		32'h0000E742: begin
				q			<=			16'h00C8;
		end
		32'h0000E744: begin
				q			<=			16'hF06F;
		end
		32'h0000E746: begin
				q			<=			16'hEC5F;
		end
		32'h0000E748: begin
				q			<=			16'h9713;
		end
		32'h0000E74A: begin
				q			<=			16'h0027;
		end
		32'h0000E74C: begin
				q			<=			16'h0613;
		end
		32'h0000E74E: begin
				q			<=			16'h0301;
		end
		32'h0000E750: begin
				q			<=			16'h0733;
		end
		32'h0000E752: begin
				q			<=			16'h00E6;
		end
		32'h0000E754: begin
				q			<=			16'h2023;
		end
		32'h0000E756: begin
				q			<=			16'h0007;
		end
		32'h0000E758: begin
				q			<=			16'h8793;
		end
		32'h0000E75A: begin
				q			<=			16'hFFF7;
		end
		32'h0000E75C: begin
				q			<=			16'hF06F;
		end
		32'h0000E75E: begin
				q			<=			16'hF4DF;
		end
		32'h0000E760: begin
				q			<=			16'h1693;
		end
		32'h0000E762: begin
				q			<=			16'h0027;
		end
		32'h0000E764: begin
				q			<=			16'h0613;
		end
		32'h0000E766: begin
				q			<=			16'h0301;
		end
		32'h0000E768: begin
				q			<=			16'h06B3;
		end
		32'h0000E76A: begin
				q			<=			16'h00D6;
		end
		32'h0000E76C: begin
				q			<=			16'hA683;
		end
		32'h0000E76E: begin
				q			<=			16'h0006;
		end
		32'h0000E770: begin
				q			<=			16'h0713;
		end
		32'h0000E772: begin
				q			<=			16'h0017;
		end
		32'h0000E774: begin
				q			<=			16'h6533;
		end
		32'h0000E776: begin
				q			<=			16'h00D5;
		end
		32'h0000E778: begin
				q			<=			16'hF06F;
		end
		32'h0000E77A: begin
				q			<=			16'hF55F;
		end
		32'h0000E77C: begin
				q			<=			16'h0633;
		end
		32'h0000E77E: begin
				q			<=			16'h0067;
		end
		32'h0000E780: begin
				q			<=			16'h2603;
		end
		32'h0000E782: begin
				q			<=			16'h0006;
		end
		32'h0000E784: begin
				q			<=			16'h0413;
		end
		32'h0000E786: begin
				q			<=			16'h0014;
		end
		32'h0000E788: begin
				q			<=			16'h0713;
		end
		32'h0000E78A: begin
				q			<=			16'h0047;
		end
		32'h0000E78C: begin
				q			<=			16'h2E23;
		end
		32'h0000E78E: begin
				q			<=			16'hFEC7;
		end
		32'h0000E790: begin
				q			<=			16'hF06F;
		end
		32'h0000E792: begin
				q			<=			16'hF61F;
		end
		32'h0000E794: begin
				q			<=			16'h1713;
		end
		32'h0000E796: begin
				q			<=			16'h0027;
		end
		32'h0000E798: begin
				q			<=			16'h0693;
		end
		32'h0000E79A: begin
				q			<=			16'h0401;
		end
		32'h0000E79C: begin
				q			<=			16'h8733;
		end
		32'h0000E79E: begin
				q			<=			16'h00E6;
		end
		32'h0000E7A0: begin
				q			<=			16'h2703;
		end
		32'h0000E7A2: begin
				q			<=			16'hFF07;
		end
		32'h0000E7A4: begin
				q			<=			16'h0613;
		end
		32'h0000E7A6: begin
				q			<=			16'h0200;
		end
		32'h0000E7A8: begin
				q			<=			16'h0633;
		end
		32'h0000E7AA: begin
				q			<=			16'h4086;
		end
		32'h0000E7AC: begin
				q			<=			16'h1733;
		end
		32'h0000E7AE: begin
				q			<=			16'h00C7;
		end
		32'h0000E7B0: begin
				q			<=			16'h6533;
		end
		32'h0000E7B2: begin
				q			<=			16'h00E5;
		end
		32'h0000E7B4: begin
				q			<=			16'h0713;
		end
		32'h0000E7B6: begin
				q			<=			16'h0030;
		end
		32'h0000E7B8: begin
				q			<=			16'h0593;
		end
		32'h0000E7BA: begin
				q			<=			16'h0301;
		end
		32'h0000E7BC: begin
				q			<=			16'h0813;
		end
		32'h0000E7BE: begin
				q			<=			16'h0000;
		end
		32'h0000E7C0: begin
				q			<=			16'h0733;
		end
		32'h0000E7C2: begin
				q			<=			16'h40F7;
		end
		32'h0000E7C4: begin
				q			<=			16'h4463;
		end
		32'h0000E7C6: begin
				q			<=			16'h02E8;
		end
		32'h0000E7C8: begin
				q			<=			16'h0693;
		end
		32'h0000E7CA: begin
				q			<=			16'h0040;
		end
		32'h0000E7CC: begin
				q			<=			16'h87B3;
		end
		32'h0000E7CE: begin
				q			<=			16'h40F6;
		end
		32'h0000E7D0: begin
				q			<=			16'h1713;
		end
		32'h0000E7D2: begin
				q			<=			16'h0027;
		end
		32'h0000E7D4: begin
				q			<=			16'h0693;
		end
		32'h0000E7D6: begin
				q			<=			16'h0401;
		end
		32'h0000E7D8: begin
				q			<=			16'h8733;
		end
		32'h0000E7DA: begin
				q			<=			16'h00E6;
		end
		32'h0000E7DC: begin
				q			<=			16'h2683;
		end
		32'h0000E7DE: begin
				q			<=			16'h03C1;
		end
		32'h0000E7E0: begin
				q			<=			16'hD433;
		end
		32'h0000E7E2: begin
				q			<=			16'h0086;
		end
		32'h0000E7E4: begin
				q			<=			16'h2823;
		end
		32'h0000E7E6: begin
				q			<=			16'hFE87;
		end
		32'h0000E7E8: begin
				q			<=			16'hF06F;
		end
		32'h0000E7EA: begin
				q			<=			16'hF15F;
		end
		32'h0000E7EC: begin
				q			<=			16'h88B3;
		end
		32'h0000E7EE: begin
				q			<=			16'h0065;
		end
		32'h0000E7F0: begin
				q			<=			16'hA683;
		end
		32'h0000E7F2: begin
				q			<=			16'h0008;
		end
		32'h0000E7F4: begin
				q			<=			16'hA883;
		end
		32'h0000E7F6: begin
				q			<=			16'h0048;
		end
		32'h0000E7F8: begin
				q			<=			16'h0813;
		end
		32'h0000E7FA: begin
				q			<=			16'h0018;
		end
		32'h0000E7FC: begin
				q			<=			16'hD6B3;
		end
		32'h0000E7FE: begin
				q			<=			16'h0086;
		end
		32'h0000E800: begin
				q			<=			16'h98B3;
		end
		32'h0000E802: begin
				q			<=			16'h00C8;
		end
		32'h0000E804: begin
				q			<=			16'hE6B3;
		end
		32'h0000E806: begin
				q			<=			16'h0116;
		end
		32'h0000E808: begin
				q			<=			16'hA023;
		end
		32'h0000E80A: begin
				q			<=			16'h00D5;
		end
		32'h0000E80C: begin
				q			<=			16'h8593;
		end
		32'h0000E80E: begin
				q			<=			16'h0045;
		end
		32'h0000E810: begin
				q			<=			16'hF06F;
		end
		32'h0000E812: begin
				q			<=			16'hFB5F;
		end
		32'h0000E814: begin
				q			<=			16'h9713;
		end
		32'h0000E816: begin
				q			<=			16'h0027;
		end
		32'h0000E818: begin
				q			<=			16'h0613;
		end
		32'h0000E81A: begin
				q			<=			16'h0301;
		end
		32'h0000E81C: begin
				q			<=			16'h0733;
		end
		32'h0000E81E: begin
				q			<=			16'h00E6;
		end
		32'h0000E820: begin
				q			<=			16'h2023;
		end
		32'h0000E822: begin
				q			<=			16'h0007;
		end
		32'h0000E824: begin
				q			<=			16'h8793;
		end
		32'h0000E826: begin
				q			<=			16'h0017;
		end
		32'h0000E828: begin
				q			<=			16'hF06F;
		end
		32'h0000E82A: begin
				q			<=			16'hED9F;
		end
		32'h0000E82C: begin
				q			<=			16'h2783;
		end
		32'h0000E82E: begin
				q			<=			16'h03C1;
		end
		32'h0000E830: begin
				q			<=			16'h0737;
		end
		32'h0000E832: begin
				q			<=			16'hFFF8;
		end
		32'h0000E834: begin
				q			<=			16'h0713;
		end
		32'h0000E836: begin
				q			<=			16'hFFF7;
		end
		32'h0000E838: begin
				q			<=			16'h0433;
		end
		32'h0000E83A: begin
				q			<=			16'h40A4;
		end
		32'h0000E83C: begin
				q			<=			16'hF7B3;
		end
		32'h0000E83E: begin
				q			<=			16'h00E7;
		end
		32'h0000E840: begin
				q			<=			16'hE06F;
		end
		32'h0000E842: begin
				q			<=			16'hE19F;
		end
		32'h0000E844: begin
				q			<=			16'h2E23;
		end
		32'h0000E846: begin
				q			<=			16'h0201;
		end
		32'h0000E848: begin
				q			<=			16'h2C23;
		end
		32'h0000E84A: begin
				q			<=			16'h0201;
		end
		32'h0000E84C: begin
				q			<=			16'h2A23;
		end
		32'h0000E84E: begin
				q			<=			16'h0201;
		end
		32'h0000E850: begin
				q			<=			16'h2823;
		end
		32'h0000E852: begin
				q			<=			16'h0201;
		end
		32'h0000E854: begin
				q			<=			16'hF06F;
		end
		32'h0000E856: begin
				q			<=			16'h854F;
		end
		32'h0000E858: begin
				q			<=			16'h0000;
		end
		32'h0000E85A: begin
				q			<=			16'h0000;
		end
		32'h0000E85C: begin
				q			<=			16'h2703;
		end
		32'h0000E85E: begin
				q			<=			16'h0045;
		end
		32'h0000E860: begin
				q			<=			16'h2783;
		end
		32'h0000E862: begin
				q			<=			16'h0085;
		end
		32'h0000E864: begin
				q			<=			16'h2603;
		end
		32'h0000E866: begin
				q			<=			16'h00C5;
		end
		32'h0000E868: begin
				q			<=			16'h2683;
		end
		32'h0000E86A: begin
				q			<=			16'h0005;
		end
		32'h0000E86C: begin
				q			<=			16'h0113;
		end
		32'h0000E86E: begin
				q			<=			16'hFE01;
		end
		32'h0000E870: begin
				q			<=			16'h2223;
		end
		32'h0000E872: begin
				q			<=			16'h00E1;
		end
		32'h0000E874: begin
				q			<=			16'h2423;
		end
		32'h0000E876: begin
				q			<=			16'h00F1;
		end
		32'h0000E878: begin
				q			<=			16'h2A23;
		end
		32'h0000E87A: begin
				q			<=			16'h00E1;
		end
		32'h0000E87C: begin
				q			<=			16'h2C23;
		end
		32'h0000E87E: begin
				q			<=			16'h00F1;
		end
		32'h0000E880: begin
				q			<=			16'h4737;
		end
		32'h0000E882: begin
				q			<=			16'h0000;
		end
		32'h0000E884: begin
				q			<=			16'h1793;
		end
		32'h0000E886: begin
				q			<=			16'h0016;
		end
		32'h0000E888: begin
				q			<=			16'h2023;
		end
		32'h0000E88A: begin
				q			<=			16'h00D1;
		end
		32'h0000E88C: begin
				q			<=			16'h2823;
		end
		32'h0000E88E: begin
				q			<=			16'h00D1;
		end
		32'h0000E890: begin
				q			<=			16'h2623;
		end
		32'h0000E892: begin
				q			<=			16'h00C1;
		end
		32'h0000E894: begin
				q			<=			16'hD693;
		end
		32'h0000E896: begin
				q			<=			16'h0117;
		end
		32'h0000E898: begin
				q			<=			16'h0793;
		end
		32'h0000E89A: begin
				q			<=			16'hFFE7;
		end
		32'h0000E89C: begin
				q			<=			16'h0513;
		end
		32'h0000E89E: begin
				q			<=			16'h0000;
		end
		32'h0000E8A0: begin
				q			<=			16'hD063;
		end
		32'h0000E8A2: begin
				q			<=			16'h02D7;
		end
		32'h0000E8A4: begin
				q			<=			16'h0793;
		end
		32'h0000E8A6: begin
				q			<=			16'h01D7;
		end
		32'h0000E8A8: begin
				q			<=			16'h1593;
		end
		32'h0000E8AA: begin
				q			<=			16'h0106;
		end
		32'h0000E8AC: begin
				q			<=			16'h5613;
		end
		32'h0000E8AE: begin
				q			<=			16'h01F6;
		end
		32'h0000E8B0: begin
				q			<=			16'hDC63;
		end
		32'h0000E8B2: begin
				q			<=			16'h00D7;
		end
		32'h0000E8B4: begin
				q			<=			16'h0537;
		end
		32'h0000E8B6: begin
				q			<=			16'h8000;
		end
		32'h0000E8B8: begin
				q			<=			16'h4513;
		end
		32'h0000E8BA: begin
				q			<=			16'hFFF5;
		end
		32'h0000E8BC: begin
				q			<=			16'h0533;
		end
		32'h0000E8BE: begin
				q			<=			16'h00A6;
		end
		32'h0000E8C0: begin
				q			<=			16'h0113;
		end
		32'h0000E8C2: begin
				q			<=			16'h0201;
		end
		32'h0000E8C4: begin
				q			<=			16'h8067;
		end
		32'h0000E8C6: begin
				q			<=			16'h0000;
		end
		32'h0000E8C8: begin
				q			<=			16'h07B7;
		end
		32'h0000E8CA: begin
				q			<=			16'h0001;
		end
		32'h0000E8CC: begin
				q			<=			16'hD593;
		end
		32'h0000E8CE: begin
				q			<=			16'h0105;
		end
		32'h0000E8D0: begin
				q			<=			16'hE5B3;
		end
		32'h0000E8D2: begin
				q			<=			16'h00F5;
		end
		32'h0000E8D4: begin
				q			<=			16'h0793;
		end
		32'h0000E8D6: begin
				q			<=			16'h06F7;
		end
		32'h0000E8D8: begin
				q			<=			16'h87B3;
		end
		32'h0000E8DA: begin
				q			<=			16'h40D7;
		end
		32'h0000E8DC: begin
				q			<=			16'hD713;
		end
		32'h0000E8DE: begin
				q			<=			16'h4057;
		end
		32'h0000E8E0: begin
				q			<=			16'h2E23;
		end
		32'h0000E8E2: begin
				q			<=			16'h00B1;
		end
		32'h0000E8E4: begin
				q			<=			16'hF793;
		end
		32'h0000E8E6: begin
				q			<=			16'h01F7;
		end
		32'h0000E8E8: begin
				q			<=			16'h9263;
		end
		32'h0000E8EA: begin
				q			<=			16'h0A07;
		end
		32'h0000E8EC: begin
				q			<=			16'h0593;
		end
		32'h0000E8EE: begin
				q			<=			16'h0030;
		end
		32'h0000E8F0: begin
				q			<=			16'h0693;
		end
		32'h0000E8F2: begin
				q			<=			16'h0101;
		end
		32'h0000E8F4: begin
				q			<=			16'h1513;
		end
		32'h0000E8F6: begin
				q			<=			16'h0027;
		end
		32'h0000E8F8: begin
				q			<=			16'h85B3;
		end
		32'h0000E8FA: begin
				q			<=			16'h40E5;
		end
		32'h0000E8FC: begin
				q			<=			16'hDE63;
		end
		32'h0000E8FE: begin
				q			<=			16'h02F5;
		end
		32'h0000E900: begin
				q			<=			16'h0793;
		end
		32'h0000E902: begin
				q			<=			16'h0040;
		end
		32'h0000E904: begin
				q			<=			16'h8733;
		end
		32'h0000E906: begin
				q			<=			16'h40E7;
		end
		32'h0000E908: begin
				q			<=			16'h0693;
		end
		32'h0000E90A: begin
				q			<=			16'h0101;
		end
		32'h0000E90C: begin
				q			<=			16'h1793;
		end
		32'h0000E90E: begin
				q			<=			16'h0027;
		end
		32'h0000E910: begin
				q			<=			16'h87B3;
		end
		32'h0000E912: begin
				q			<=			16'h00F6;
		end
		32'h0000E914: begin
				q			<=			16'h0693;
		end
		32'h0000E916: begin
				q			<=			16'h0040;
		end
		32'h0000E918: begin
				q			<=			16'hA023;
		end
		32'h0000E91A: begin
				q			<=			16'h0007;
		end
		32'h0000E91C: begin
				q			<=			16'h0713;
		end
		32'h0000E91E: begin
				q			<=			16'h0017;
		end
		32'h0000E920: begin
				q			<=			16'h8793;
		end
		32'h0000E922: begin
				q			<=			16'h0047;
		end
		32'h0000E924: begin
				q			<=			16'h1AE3;
		end
		32'h0000E926: begin
				q			<=			16'hFED7;
		end
		32'h0000E928: begin
				q			<=			16'h2503;
		end
		32'h0000E92A: begin
				q			<=			16'h0101;
		end
		32'h0000E92C: begin
				q			<=			16'h0AE3;
		end
		32'h0000E92E: begin
				q			<=			16'hF806;
		end
		32'h0000E930: begin
				q			<=			16'h0533;
		end
		32'h0000E932: begin
				q			<=			16'h40A0;
		end
		32'h0000E934: begin
				q			<=			16'hF06F;
		end
		32'h0000E936: begin
				q			<=			16'hF8DF;
		end
		32'h0000E938: begin
				q			<=			16'h8833;
		end
		32'h0000E93A: begin
				q			<=			16'h00A6;
		end
		32'h0000E93C: begin
				q			<=			16'h2803;
		end
		32'h0000E93E: begin
				q			<=			16'h0008;
		end
		32'h0000E940: begin
				q			<=			16'h8793;
		end
		32'h0000E942: begin
				q			<=			16'h0017;
		end
		32'h0000E944: begin
				q			<=			16'h8693;
		end
		32'h0000E946: begin
				q			<=			16'h0046;
		end
		32'h0000E948: begin
				q			<=			16'hAE23;
		end
		32'h0000E94A: begin
				q			<=			16'hFF06;
		end
		32'h0000E94C: begin
				q			<=			16'hF06F;
		end
		32'h0000E94E: begin
				q			<=			16'hFB1F;
		end
		32'h0000E950: begin
				q			<=			16'h2683;
		end
		32'h0000E952: begin
				q			<=			16'hFF05;
		end
		32'h0000E954: begin
				q			<=			16'h2303;
		end
		32'h0000E956: begin
				q			<=			16'hFF07;
		end
		32'h0000E958: begin
				q			<=			16'h96B3;
		end
		32'h0000E95A: begin
				q			<=			16'h0116;
		end
		32'h0000E95C: begin
				q			<=			16'h5333;
		end
		32'h0000E95E: begin
				q			<=			16'h00F3;
		end
		32'h0000E960: begin
				q			<=			16'hE6B3;
		end
		32'h0000E962: begin
				q			<=			16'h0066;
		end
		32'h0000E964: begin
				q			<=			16'h2823;
		end
		32'h0000E966: begin
				q			<=			16'h00D1;
		end
		32'h0000E968: begin
				q			<=			16'h0693;
		end
		32'h0000E96A: begin
				q			<=			16'h0010;
		end
		32'h0000E96C: begin
				q			<=			16'hC2E3;
		end
		32'h0000E96E: begin
				q			<=			16'hFF06;
		end
		32'h0000E970: begin
				q			<=			16'h8713;
		end
		32'h0000E972: begin
				q			<=			16'h0016;
		end
		32'h0000E974: begin
				q			<=			16'h0513;
		end
		32'h0000E976: begin
				q			<=			16'h0201;
		end
		32'h0000E978: begin
				q			<=			16'h9693;
		end
		32'h0000E97A: begin
				q			<=			16'h0026;
		end
		32'h0000E97C: begin
				q			<=			16'h06B3;
		end
		32'h0000E97E: begin
				q			<=			16'h00D5;
		end
		32'h0000E980: begin
				q			<=			16'hD7B3;
		end
		32'h0000E982: begin
				q			<=			16'h00F5;
		end
		32'h0000E984: begin
				q			<=			16'hA823;
		end
		32'h0000E986: begin
				q			<=			16'hFEF6;
		end
		32'h0000E988: begin
				q			<=			16'hF06F;
		end
		32'h0000E98A: begin
				q			<=			16'hF81F;
		end
		32'h0000E98C: begin
				q			<=			16'h0513;
		end
		32'h0000E98E: begin
				q			<=			16'h0017;
		end
		32'h0000E990: begin
				q			<=			16'h0893;
		end
		32'h0000E992: begin
				q			<=			16'h0201;
		end
		32'h0000E994: begin
				q			<=			16'h0813;
		end
		32'h0000E996: begin
				q			<=			16'h0030;
		end
		32'h0000E998: begin
				q			<=			16'h1513;
		end
		32'h0000E99A: begin
				q			<=			16'h0025;
		end
		32'h0000E99C: begin
				q			<=			16'h0833;
		end
		32'h0000E99E: begin
				q			<=			16'h40E8;
		end
		32'h0000E9A0: begin
				q			<=			16'h8533;
		end
		32'h0000E9A2: begin
				q			<=			16'h00A8;
		end
		32'h0000E9A4: begin
				q			<=			16'h1713;
		end
		32'h0000E9A6: begin
				q			<=			16'h0027;
		end
		32'h0000E9A8: begin
				q			<=			16'h0893;
		end
		32'h0000E9AA: begin
				q			<=			16'h0200;
		end
		32'h0000E9AC: begin
				q			<=			16'h0313;
		end
		32'h0000E9AE: begin
				q			<=			16'h0201;
		end
		32'h0000E9B0: begin
				q			<=			16'h0693;
		end
		32'h0000E9B2: begin
				q			<=			16'h0000;
		end
		32'h0000E9B4: begin
				q			<=			16'h88B3;
		end
		32'h0000E9B6: begin
				q			<=			16'h40F8;
		end
		32'h0000E9B8: begin
				q			<=			16'h0733;
		end
		32'h0000E9BA: begin
				q			<=			16'h00E3;
		end
		32'h0000E9BC: begin
				q			<=			16'hF06F;
		end
		32'h0000E9BE: begin
				q			<=			16'hFB1F;
		end
		32'h0000E9C0: begin
				q			<=			16'h0000;
		end
		32'h0000E9C2: begin
				q			<=			16'h0000;
		end
		32'h0000E9C4: begin
				q			<=			16'h0113;
		end
		32'h0000E9C6: begin
				q			<=			16'hFD01;
		end
		32'h0000E9C8: begin
				q			<=			16'h2223;
		end
		32'h0000E9CA: begin
				q			<=			16'h0291;
		end
		32'h0000E9CC: begin
				q			<=			16'h2623;
		end
		32'h0000E9CE: begin
				q			<=			16'h0211;
		end
		32'h0000E9D0: begin
				q			<=			16'h2423;
		end
		32'h0000E9D2: begin
				q			<=			16'h0281;
		end
		32'h0000E9D4: begin
				q			<=			16'h2023;
		end
		32'h0000E9D6: begin
				q			<=			16'h0321;
		end
		32'h0000E9D8: begin
				q			<=			16'h0493;
		end
		32'h0000E9DA: begin
				q			<=			16'h0005;
		end
		32'h0000E9DC: begin
				q			<=			16'h8663;
		end
		32'h0000E9DE: begin
				q			<=			16'h1405;
		end
		32'h0000E9E0: begin
				q			<=			16'h8413;
		end
		32'h0000E9E2: begin
				q			<=			16'h0005;
		end
		32'h0000E9E4: begin
				q			<=			16'hD913;
		end
		32'h0000E9E6: begin
				q			<=			16'h01F5;
		end
		32'h0000E9E8: begin
				q			<=			16'hD463;
		end
		32'h0000E9EA: begin
				q			<=			16'h0005;
		end
		32'h0000E9EC: begin
				q			<=			16'h0433;
		end
		32'h0000E9EE: begin
				q			<=			16'h40B0;
		end
		32'h0000E9F0: begin
				q			<=			16'h0513;
		end
		32'h0000E9F2: begin
				q			<=			16'h0004;
		end
		32'h0000E9F4: begin
				q			<=			16'h00EF;
		end
		32'h0000E9F6: begin
				q			<=			16'h6D80;
		end
		32'h0000E9F8: begin
				q			<=			16'h0593;
		end
		32'h0000E9FA: begin
				q			<=			16'h0515;
		end
		32'h0000E9FC: begin
				q			<=			16'h4737;
		end
		32'h0000E9FE: begin
				q			<=			16'h0000;
		end
		32'h0000EA00: begin
				q			<=			16'h0713;
		end
		32'h0000EA02: begin
				q			<=			16'h01E7;
		end
		32'h0000EA04: begin
				q			<=			16'hD793;
		end
		32'h0000EA06: begin
				q			<=			16'h4055;
		end
		32'h0000EA08: begin
				q			<=			16'h2823;
		end
		32'h0000EA0A: begin
				q			<=			16'h0081;
		end
		32'h0000EA0C: begin
				q			<=			16'h2A23;
		end
		32'h0000EA0E: begin
				q			<=			16'h0001;
		end
		32'h0000EA10: begin
				q			<=			16'h2C23;
		end
		32'h0000EA12: begin
				q			<=			16'h0001;
		end
		32'h0000EA14: begin
				q			<=			16'h2E23;
		end
		32'h0000EA16: begin
				q			<=			16'h0001;
		end
		32'h0000EA18: begin
				q			<=			16'hF593;
		end
		32'h0000EA1A: begin
				q			<=			16'h01F5;
		end
		32'h0000EA1C: begin
				q			<=			16'h0733;
		end
		32'h0000EA1E: begin
				q			<=			16'h40A7;
		end
		32'h0000EA20: begin
				q			<=			16'h8C63;
		end
		32'h0000EA22: begin
				q			<=			16'h0205;
		end
		32'h0000EA24: begin
				q			<=			16'h0693;
		end
		32'h0000EA26: begin
				q			<=			16'h0020;
		end
		32'h0000EA28: begin
				q			<=			16'h9C63;
		end
		32'h0000EA2A: begin
				q			<=			16'h0ED7;
		end
		32'h0000EA2C: begin
				q			<=			16'h0693;
		end
		32'h0000EA2E: begin
				q			<=			16'h0200;
		end
		32'h0000EA30: begin
				q			<=			16'h86B3;
		end
		32'h0000EA32: begin
				q			<=			16'h40B6;
		end
		32'h0000EA34: begin
				q			<=			16'h56B3;
		end
		32'h0000EA36: begin
				q			<=			16'h00D4;
		end
		32'h0000EA38: begin
				q			<=			16'h2E23;
		end
		32'h0000EA3A: begin
				q			<=			16'h00D1;
		end
		32'h0000EA3C: begin
				q			<=			16'h8693;
		end
		32'h0000EA3E: begin
				q			<=			16'hFFF7;
		end
		32'h0000EA40: begin
				q			<=			16'h0613;
		end
		32'h0000EA42: begin
				q			<=			16'h0201;
		end
		32'h0000EA44: begin
				q			<=			16'h9793;
		end
		32'h0000EA46: begin
				q			<=			16'h0027;
		end
		32'h0000EA48: begin
				q			<=			16'h07B3;
		end
		32'h0000EA4A: begin
				q			<=			16'h00F6;
		end
		32'h0000EA4C: begin
				q			<=			16'h1433;
		end
		32'h0000EA4E: begin
				q			<=			16'h00B4;
		end
		32'h0000EA50: begin
				q			<=			16'hA823;
		end
		32'h0000EA52: begin
				q			<=			16'hFE87;
		end
		32'h0000EA54: begin
				q			<=			16'h006F;
		end
		32'h0000EA56: begin
				q			<=			16'h0340;
		end
		32'h0000EA58: begin
				q			<=			16'h0693;
		end
		32'h0000EA5A: begin
				q			<=			16'h0030;
		end
		32'h0000EA5C: begin
				q			<=			16'h86B3;
		end
		32'h0000EA5E: begin
				q			<=			16'h40F6;
		end
		32'h0000EA60: begin
				q			<=			16'h0613;
		end
		32'h0000EA62: begin
				q			<=			16'h0201;
		end
		32'h0000EA64: begin
				q			<=			16'h9693;
		end
		32'h0000EA66: begin
				q			<=			16'h0026;
		end
		32'h0000EA68: begin
				q			<=			16'h06B3;
		end
		32'h0000EA6A: begin
				q			<=			16'h00D6;
		end
		32'h0000EA6C: begin
				q			<=			16'hA683;
		end
		32'h0000EA6E: begin
				q			<=			16'hFF06;
		end
		32'h0000EA70: begin
				q			<=			16'h0613;
		end
		32'h0000EA72: begin
				q			<=			16'h0020;
		end
		32'h0000EA74: begin
				q			<=			16'h2E23;
		end
		32'h0000EA76: begin
				q			<=			16'h00D1;
		end
		32'h0000EA78: begin
				q			<=			16'h0693;
		end
		32'h0000EA7A: begin
				q			<=			16'h0020;
		end
		32'h0000EA7C: begin
				q			<=			16'h9663;
		end
		32'h0000EA7E: begin
				q			<=			16'h00C7;
		end
		32'h0000EA80: begin
				q			<=			16'h2C23;
		end
		32'h0000EA82: begin
				q			<=			16'h0081;
		end
		32'h0000EA84: begin
				q			<=			16'h0693;
		end
		32'h0000EA86: begin
				q			<=			16'h0010;
		end
		32'h0000EA88: begin
				q			<=			16'h0793;
		end
		32'h0000EA8A: begin
				q			<=			16'h0101;
		end
		32'h0000EA8C: begin
				q			<=			16'h9613;
		end
		32'h0000EA8E: begin
				q			<=			16'h0026;
		end
		32'h0000EA90: begin
				q			<=			16'h8633;
		end
		32'h0000EA92: begin
				q			<=			16'h00C7;
		end
		32'h0000EA94: begin
				q			<=			16'h0793;
		end
		32'h0000EA96: begin
				q			<=			16'hFFF0;
		end
		32'h0000EA98: begin
				q			<=			16'h2023;
		end
		32'h0000EA9A: begin
				q			<=			16'h0006;
		end
		32'h0000EA9C: begin
				q			<=			16'h8693;
		end
		32'h0000EA9E: begin
				q			<=			16'hFFF6;
		end
		32'h0000EAA0: begin
				q			<=			16'h0613;
		end
		32'h0000EAA2: begin
				q			<=			16'hFFC6;
		end
		32'h0000EAA4: begin
				q			<=			16'h9AE3;
		end
		32'h0000EAA6: begin
				q			<=			16'hFEF6;
		end
		32'h0000EAA8: begin
				q			<=			16'h86B7;
		end
		32'h0000EAAA: begin
				q			<=			16'h0000;
		end
		32'h0000EAAC: begin
				q			<=			16'h2783;
		end
		32'h0000EAAE: begin
				q			<=			16'h01C1;
		end
		32'h0000EAB0: begin
				q			<=			16'h8693;
		end
		32'h0000EAB2: begin
				q			<=			16'hFFF6;
		end
		32'h0000EAB4: begin
				q			<=			16'h76B3;
		end
		32'h0000EAB6: begin
				q			<=			16'h00D7;
		end
		32'h0000EAB8: begin
				q			<=			16'h5703;
		end
		32'h0000EABA: begin
				q			<=			16'h00E1;
		end
		32'h0000EABC: begin
				q			<=			16'h1623;
		end
		32'h0000EABE: begin
				q			<=			16'h00F1;
		end
		32'h0000EAC0: begin
				q			<=			16'h87B7;
		end
		32'h0000EAC2: begin
				q			<=			16'hFFFF;
		end
		32'h0000EAC4: begin
				q			<=			16'h7733;
		end
		32'h0000EAC6: begin
				q			<=			16'h00F7;
		end
		32'h0000EAC8: begin
				q			<=			16'h6733;
		end
		32'h0000EACA: begin
				q			<=			16'h00D7;
		end
		32'h0000EACC: begin
				q			<=			16'h5793;
		end
		32'h0000EACE: begin
				q			<=			16'h0087;
		end
		32'h0000EAD0: begin
				q			<=			16'h1723;
		end
		32'h0000EAD2: begin
				q			<=			16'h00E1;
		end
		32'h0000EAD4: begin
				q			<=			16'hF793;
		end
		32'h0000EAD6: begin
				q			<=			16'h07F7;
		end
		32'h0000EAD8: begin
				q			<=			16'h1713;
		end
		32'h0000EADA: begin
				q			<=			16'h0079;
		end
		32'h0000EADC: begin
				q			<=			16'hE7B3;
		end
		32'h0000EADE: begin
				q			<=			16'h00E7;
		end
		32'h0000EAE0: begin
				q			<=			16'h07A3;
		end
		32'h0000EAE2: begin
				q			<=			16'h00F1;
		end
		32'h0000EAE4: begin
				q			<=			16'h2783;
		end
		32'h0000EAE6: begin
				q			<=			16'h0101;
		end
		32'h0000EAE8: begin
				q			<=			16'h2083;
		end
		32'h0000EAEA: begin
				q			<=			16'h02C1;
		end
		32'h0000EAEC: begin
				q			<=			16'h2403;
		end
		32'h0000EAEE: begin
				q			<=			16'h0281;
		end
		32'h0000EAF0: begin
				q			<=			16'hA023;
		end
		32'h0000EAF2: begin
				q			<=			16'h00F4;
		end
		32'h0000EAF4: begin
				q			<=			16'h2783;
		end
		32'h0000EAF6: begin
				q			<=			16'h0141;
		end
		32'h0000EAF8: begin
				q			<=			16'h8513;
		end
		32'h0000EAFA: begin
				q			<=			16'h0004;
		end
		32'h0000EAFC: begin
				q			<=			16'h2903;
		end
		32'h0000EAFE: begin
				q			<=			16'h0201;
		end
		32'h0000EB00: begin
				q			<=			16'hA223;
		end
		32'h0000EB02: begin
				q			<=			16'h00F4;
		end
		32'h0000EB04: begin
				q			<=			16'h2783;
		end
		32'h0000EB06: begin
				q			<=			16'h0181;
		end
		32'h0000EB08: begin
				q			<=			16'hA423;
		end
		32'h0000EB0A: begin
				q			<=			16'h00F4;
		end
		32'h0000EB0C: begin
				q			<=			16'h2783;
		end
		32'h0000EB0E: begin
				q			<=			16'h00C1;
		end
		32'h0000EB10: begin
				q			<=			16'hA623;
		end
		32'h0000EB12: begin
				q			<=			16'h00F4;
		end
		32'h0000EB14: begin
				q			<=			16'h2483;
		end
		32'h0000EB16: begin
				q			<=			16'h0241;
		end
		32'h0000EB18: begin
				q			<=			16'h0113;
		end
		32'h0000EB1A: begin
				q			<=			16'h0301;
		end
		32'h0000EB1C: begin
				q			<=			16'h8067;
		end
		32'h0000EB1E: begin
				q			<=			16'h0000;
		end
		32'h0000EB20: begin
				q			<=			16'h0793;
		end
		32'h0000EB22: begin
				q			<=			16'h0030;
		end
		32'h0000EB24: begin
				q			<=			16'hF06F;
		end
		32'h0000EB26: begin
				q			<=			16'hF19F;
		end
		32'h0000EB28: begin
				q			<=			16'h2E23;
		end
		32'h0000EB2A: begin
				q			<=			16'h0001;
		end
		32'h0000EB2C: begin
				q			<=			16'h2C23;
		end
		32'h0000EB2E: begin
				q			<=			16'h0001;
		end
		32'h0000EB30: begin
				q			<=			16'h2A23;
		end
		32'h0000EB32: begin
				q			<=			16'h0001;
		end
		32'h0000EB34: begin
				q			<=			16'h2823;
		end
		32'h0000EB36: begin
				q			<=			16'h0001;
		end
		32'h0000EB38: begin
				q			<=			16'h0713;
		end
		32'h0000EB3A: begin
				q			<=			16'h0000;
		end
		32'h0000EB3C: begin
				q			<=			16'h0913;
		end
		32'h0000EB3E: begin
				q			<=			16'h0000;
		end
		32'h0000EB40: begin
				q			<=			16'hF06F;
		end
		32'h0000EB42: begin
				q			<=			16'hF69F;
		end
		32'h0000EB44: begin
				q			<=			16'h0000;
		end
		32'h0000EB46: begin
				q			<=			16'h0000;
		end
		32'h0000EB48: begin
				q			<=			16'h5793;
		end
		32'h0000EB4A: begin
				q			<=			16'h0146;
		end
		32'h0000EB4C: begin
				q			<=			16'h0737;
		end
		32'h0000EB4E: begin
				q			<=			16'h0010;
		end
		32'h0000EB50: begin
				q			<=			16'h0713;
		end
		32'h0000EB52: begin
				q			<=			16'hFFF7;
		end
		32'h0000EB54: begin
				q			<=			16'hF793;
		end
		32'h0000EB56: begin
				q			<=			16'h7FF7;
		end
		32'h0000EB58: begin
				q			<=			16'h0113;
		end
		32'h0000EB5A: begin
				q			<=			16'hFD01;
		end
		32'h0000EB5C: begin
				q			<=			16'h7733;
		end
		32'h0000EB5E: begin
				q			<=			16'h00C7;
		end
		32'h0000EB60: begin
				q			<=			16'h8693;
		end
		32'h0000EB62: begin
				q			<=			16'h0017;
		end
		32'h0000EB64: begin
				q			<=			16'h2423;
		end
		32'h0000EB66: begin
				q			<=			16'h0281;
		end
		32'h0000EB68: begin
				q			<=			16'h2223;
		end
		32'h0000EB6A: begin
				q			<=			16'h0291;
		end
		32'h0000EB6C: begin
				q			<=			16'h5413;
		end
		32'h0000EB6E: begin
				q			<=			16'h01F6;
		end
		32'h0000EB70: begin
				q			<=			16'h2623;
		end
		32'h0000EB72: begin
				q			<=			16'h0211;
		end
		32'h0000EB74: begin
				q			<=			16'h2823;
		end
		32'h0000EB76: begin
				q			<=			16'h00B1;
		end
		32'h0000EB78: begin
				q			<=			16'h2A23;
		end
		32'h0000EB7A: begin
				q			<=			16'h00E1;
		end
		32'h0000EB7C: begin
				q			<=			16'h2E23;
		end
		32'h0000EB7E: begin
				q			<=			16'h0001;
		end
		32'h0000EB80: begin
				q			<=			16'h2C23;
		end
		32'h0000EB82: begin
				q			<=			16'h0001;
		end
		32'h0000EB84: begin
				q			<=			16'hF693;
		end
		32'h0000EB86: begin
				q			<=			16'h7FF6;
		end
		32'h0000EB88: begin
				q			<=			16'h0613;
		end
		32'h0000EB8A: begin
				q			<=			16'h0010;
		end
		32'h0000EB8C: begin
				q			<=			16'h0493;
		end
		32'h0000EB8E: begin
				q			<=			16'h0005;
		end
		32'h0000EB90: begin
				q			<=			16'h5463;
		end
		32'h0000EB92: begin
				q			<=			16'h0AD6;
		end
		32'h0000EB94: begin
				q			<=			16'h46B7;
		end
		32'h0000EB96: begin
				q			<=			16'h0000;
		end
		32'h0000EB98: begin
				q			<=			16'h8693;
		end
		32'h0000EB9A: begin
				q			<=			16'hC006;
		end
		32'h0000EB9C: begin
				q			<=			16'hD513;
		end
		32'h0000EB9E: begin
				q			<=			16'h0045;
		end
		32'h0000EBA0: begin
				q			<=			16'h87B3;
		end
		32'h0000EBA2: begin
				q			<=			16'h00D7;
		end
		32'h0000EBA4: begin
				q			<=			16'h5693;
		end
		32'h0000EBA6: begin
				q			<=			16'h0047;
		end
		32'h0000EBA8: begin
				q			<=			16'h1713;
		end
		32'h0000EBAA: begin
				q			<=			16'h01C7;
		end
		32'h0000EBAC: begin
				q			<=			16'h6733;
		end
		32'h0000EBAE: begin
				q			<=			16'h00A7;
		end
		32'h0000EBB0: begin
				q			<=			16'h9593;
		end
		32'h0000EBB2: begin
				q			<=			16'h01C5;
		end
		32'h0000EBB4: begin
				q			<=			16'h2E23;
		end
		32'h0000EBB6: begin
				q			<=			16'h00D1;
		end
		32'h0000EBB8: begin
				q			<=			16'h2C23;
		end
		32'h0000EBBA: begin
				q			<=			16'h00E1;
		end
		32'h0000EBBC: begin
				q			<=			16'h2A23;
		end
		32'h0000EBBE: begin
				q			<=			16'h00B1;
		end
		32'h0000EBC0: begin
				q			<=			16'h2823;
		end
		32'h0000EBC2: begin
				q			<=			16'h0001;
		end
		32'h0000EBC4: begin
				q			<=			16'h8537;
		end
		32'h0000EBC6: begin
				q			<=			16'h0000;
		end
		32'h0000EBC8: begin
				q			<=			16'h2703;
		end
		32'h0000EBCA: begin
				q			<=			16'h01C1;
		end
		32'h0000EBCC: begin
				q			<=			16'h0513;
		end
		32'h0000EBCE: begin
				q			<=			16'hFFF5;
		end
		32'h0000EBD0: begin
				q			<=			16'hF7B3;
		end
		32'h0000EBD2: begin
				q			<=			16'h00A7;
		end
		32'h0000EBD4: begin
				q			<=			16'h5503;
		end
		32'h0000EBD6: begin
				q			<=			16'h00E1;
		end
		32'h0000EBD8: begin
				q			<=			16'h1623;
		end
		32'h0000EBDA: begin
				q			<=			16'h00E1;
		end
		32'h0000EBDC: begin
				q			<=			16'h8737;
		end
		32'h0000EBDE: begin
				q			<=			16'hFFFF;
		end
		32'h0000EBE0: begin
				q			<=			16'h7533;
		end
		32'h0000EBE2: begin
				q			<=			16'h00E5;
		end
		32'h0000EBE4: begin
				q			<=			16'h67B3;
		end
		32'h0000EBE6: begin
				q			<=			16'h00F5;
		end
		32'h0000EBE8: begin
				q			<=			16'h1723;
		end
		32'h0000EBEA: begin
				q			<=			16'h00F1;
		end
		32'h0000EBEC: begin
				q			<=			16'hD713;
		end
		32'h0000EBEE: begin
				q			<=			16'h0087;
		end
		32'h0000EBF0: begin
				q			<=			16'h2783;
		end
		32'h0000EBF2: begin
				q			<=			16'h0101;
		end
		32'h0000EBF4: begin
				q			<=			16'h1613;
		end
		32'h0000EBF6: begin
				q			<=			16'h0074;
		end
		32'h0000EBF8: begin
				q			<=			16'h7413;
		end
		32'h0000EBFA: begin
				q			<=			16'h07F7;
		end
		32'h0000EBFC: begin
				q			<=			16'hA023;
		end
		32'h0000EBFE: begin
				q			<=			16'h00F4;
		end
		32'h0000EC00: begin
				q			<=			16'h2783;
		end
		32'h0000EC02: begin
				q			<=			16'h0141;
		end
		32'h0000EC04: begin
				q			<=			16'h6433;
		end
		32'h0000EC06: begin
				q			<=			16'h00C4;
		end
		32'h0000EC08: begin
				q			<=			16'h07A3;
		end
		32'h0000EC0A: begin
				q			<=			16'h0081;
		end
		32'h0000EC0C: begin
				q			<=			16'hA223;
		end
		32'h0000EC0E: begin
				q			<=			16'h00F4;
		end
		32'h0000EC10: begin
				q			<=			16'h2783;
		end
		32'h0000EC12: begin
				q			<=			16'h0181;
		end
		32'h0000EC14: begin
				q			<=			16'h2083;
		end
		32'h0000EC16: begin
				q			<=			16'h02C1;
		end
		32'h0000EC18: begin
				q			<=			16'h2403;
		end
		32'h0000EC1A: begin
				q			<=			16'h0281;
		end
		32'h0000EC1C: begin
				q			<=			16'hA423;
		end
		32'h0000EC1E: begin
				q			<=			16'h00F4;
		end
		32'h0000EC20: begin
				q			<=			16'h2783;
		end
		32'h0000EC22: begin
				q			<=			16'h00C1;
		end
		32'h0000EC24: begin
				q			<=			16'h8513;
		end
		32'h0000EC26: begin
				q			<=			16'h0004;
		end
		32'h0000EC28: begin
				q			<=			16'hA623;
		end
		32'h0000EC2A: begin
				q			<=			16'h00F4;
		end
		32'h0000EC2C: begin
				q			<=			16'h2483;
		end
		32'h0000EC2E: begin
				q			<=			16'h0241;
		end
		32'h0000EC30: begin
				q			<=			16'h0113;
		end
		32'h0000EC32: begin
				q			<=			16'h0301;
		end
		32'h0000EC34: begin
				q			<=			16'h8067;
		end
		32'h0000EC36: begin
				q			<=			16'h0000;
		end
		32'h0000EC38: begin
				q			<=			16'h6533;
		end
		32'h0000EC3A: begin
				q			<=			16'h00B7;
		end
		32'h0000EC3C: begin
				q			<=			16'h9A63;
		end
		32'h0000EC3E: begin
				q			<=			16'h0E07;
		end
		32'h0000EC40: begin
				q			<=			16'h02E3;
		end
		32'h0000EC42: begin
				q			<=			16'hF805;
		end
		32'h0000EC44: begin
				q			<=			16'h0063;
		end
		32'h0000EC46: begin
				q			<=			16'h0607;
		end
		32'h0000EC48: begin
				q			<=			16'h0513;
		end
		32'h0000EC4A: begin
				q			<=			16'h0007;
		end
		32'h0000EC4C: begin
				q			<=			16'h00EF;
		end
		32'h0000EC4E: begin
				q			<=			16'h4800;
		end
		32'h0000EC50: begin
				q			<=			16'h0693;
		end
		32'h0000EC52: begin
				q			<=			16'h0315;
		end
		32'h0000EC54: begin
				q			<=			16'hD713;
		end
		32'h0000EC56: begin
				q			<=			16'h4056;
		end
		32'h0000EC58: begin
				q			<=			16'hF693;
		end
		32'h0000EC5A: begin
				q			<=			16'h01F6;
		end
		32'h0000EC5C: begin
				q			<=			16'h8A63;
		end
		32'h0000EC5E: begin
				q			<=			16'h0406;
		end
		32'h0000EC60: begin
				q			<=			16'h0613;
		end
		32'h0000EC62: begin
				q			<=			16'hFFC0;
		end
		32'h0000EC64: begin
				q			<=			16'h0633;
		end
		32'h0000EC66: begin
				q			<=			16'h02C7;
		end
		32'h0000EC68: begin
				q			<=			16'h0813;
		end
		32'h0000EC6A: begin
				q			<=			16'h0200;
		end
		32'h0000EC6C: begin
				q			<=			16'h0793;
		end
		32'h0000EC6E: begin
				q			<=			16'h0101;
		end
		32'h0000EC70: begin
				q			<=			16'h0313;
		end
		32'h0000EC72: begin
				q			<=			16'hFF00;
		end
		32'h0000EC74: begin
				q			<=			16'h0833;
		end
		32'h0000EC76: begin
				q			<=			16'h40D8;
		end
		32'h0000EC78: begin
				q			<=			16'h0613;
		end
		32'h0000EC7A: begin
				q			<=			16'hFFC6;
		end
		32'h0000EC7C: begin
				q			<=			16'h8793;
		end
		32'h0000EC7E: begin
				q			<=			16'hFFC7;
		end
		32'h0000EC80: begin
				q			<=			16'h1663;
		end
		32'h0000EC82: begin
				q			<=			16'h0866;
		end
		32'h0000EC84: begin
				q			<=			16'h0793;
		end
		32'h0000EC86: begin
				q			<=			16'h0201;
		end
		32'h0000EC88: begin
				q			<=			16'h0613;
		end
		32'h0000EC8A: begin
				q			<=			16'hFFF7;
		end
		32'h0000EC8C: begin
				q			<=			16'h1713;
		end
		32'h0000EC8E: begin
				q			<=			16'h0027;
		end
		32'h0000EC90: begin
				q			<=			16'h8733;
		end
		32'h0000EC92: begin
				q			<=			16'h00E7;
		end
		32'h0000EC94: begin
				q			<=			16'h2783;
		end
		32'h0000EC96: begin
				q			<=			16'h0101;
		end
		32'h0000EC98: begin
				q			<=			16'h96B3;
		end
		32'h0000EC9A: begin
				q			<=			16'h00D7;
		end
		32'h0000EC9C: begin
				q			<=			16'h2823;
		end
		32'h0000EC9E: begin
				q			<=			16'hFED7;
		end
		32'h0000ECA0: begin
				q			<=			16'h006F;
		end
		32'h0000ECA2: begin
				q			<=			16'h03C0;
		end
		32'h0000ECA4: begin
				q			<=			16'h00EF;
		end
		32'h0000ECA6: begin
				q			<=			16'h4280;
		end
		32'h0000ECA8: begin
				q			<=			16'h0513;
		end
		32'h0000ECAA: begin
				q			<=			16'h0205;
		end
		32'h0000ECAC: begin
				q			<=			16'hF06F;
		end
		32'h0000ECAE: begin
				q			<=			16'hFA5F;
		end
		32'h0000ECB0: begin
				q			<=			16'h0613;
		end
		32'h0000ECB2: begin
				q			<=			16'hFFC0;
		end
		32'h0000ECB4: begin
				q			<=			16'h0633;
		end
		32'h0000ECB6: begin
				q			<=			16'h02C7;
		end
		32'h0000ECB8: begin
				q			<=			16'h0693;
		end
		32'h0000ECBA: begin
				q			<=			16'h0101;
		end
		32'h0000ECBC: begin
				q			<=			16'h0793;
		end
		32'h0000ECBE: begin
				q			<=			16'h0030;
		end
		32'h0000ECC0: begin
				q			<=			16'h85B3;
		end
		32'h0000ECC2: begin
				q			<=			16'h00C6;
		end
		32'h0000ECC4: begin
				q			<=			16'hA583;
		end
		32'h0000ECC6: begin
				q			<=			16'h00C5;
		end
		32'h0000ECC8: begin
				q			<=			16'h8793;
		end
		32'h0000ECCA: begin
				q			<=			16'hFFF7;
		end
		32'h0000ECCC: begin
				q			<=			16'h8693;
		end
		32'h0000ECCE: begin
				q			<=			16'hFFC6;
		end
		32'h0000ECD0: begin
				q			<=			16'hA823;
		end
		32'h0000ECD2: begin
				q			<=			16'h00B6;
		end
		32'h0000ECD4: begin
				q			<=			16'hD6E3;
		end
		32'h0000ECD6: begin
				q			<=			16'hFEE7;
		end
		32'h0000ECD8: begin
				q			<=			16'h0613;
		end
		32'h0000ECDA: begin
				q			<=			16'hFFF7;
		end
		32'h0000ECDC: begin
				q			<=			16'h0793;
		end
		32'h0000ECDE: begin
				q			<=			16'h0101;
		end
		32'h0000ECE0: begin
				q			<=			16'h1713;
		end
		32'h0000ECE2: begin
				q			<=			16'h0026;
		end
		32'h0000ECE4: begin
				q			<=			16'h8733;
		end
		32'h0000ECE6: begin
				q			<=			16'h00E7;
		end
		32'h0000ECE8: begin
				q			<=			16'h0793;
		end
		32'h0000ECEA: begin
				q			<=			16'hFFF0;
		end
		32'h0000ECEC: begin
				q			<=			16'h2023;
		end
		32'h0000ECEE: begin
				q			<=			16'h0007;
		end
		32'h0000ECF0: begin
				q			<=			16'h0613;
		end
		32'h0000ECF2: begin
				q			<=			16'hFFF6;
		end
		32'h0000ECF4: begin
				q			<=			16'h0713;
		end
		32'h0000ECF6: begin
				q			<=			16'hFFC7;
		end
		32'h0000ECF8: begin
				q			<=			16'h1AE3;
		end
		32'h0000ECFA: begin
				q			<=			16'hFEF6;
		end
		32'h0000ECFC: begin
				q			<=			16'h47B7;
		end
		32'h0000ECFE: begin
				q			<=			16'h0000;
		end
		32'h0000ED00: begin
				q			<=			16'h8793;
		end
		32'h0000ED02: begin
				q			<=			16'hC0C7;
		end
		32'h0000ED04: begin
				q			<=			16'h87B3;
		end
		32'h0000ED06: begin
				q			<=			16'h40A7;
		end
		32'h0000ED08: begin
				q			<=			16'hF06F;
		end
		32'h0000ED0A: begin
				q			<=			16'hEBDF;
		end
		32'h0000ED0C: begin
				q			<=			16'h0593;
		end
		32'h0000ED0E: begin
				q			<=			16'h0101;
		end
		32'h0000ED10: begin
				q			<=			16'h88B3;
		end
		32'h0000ED12: begin
				q			<=			16'h00C5;
		end
		32'h0000ED14: begin
				q			<=			16'hA583;
		end
		32'h0000ED16: begin
				q			<=			16'h00C8;
		end
		32'h0000ED18: begin
				q			<=			16'hA883;
		end
		32'h0000ED1A: begin
				q			<=			16'h0108;
		end
		32'h0000ED1C: begin
				q			<=			16'hD5B3;
		end
		32'h0000ED1E: begin
				q			<=			16'h0105;
		end
		32'h0000ED20: begin
				q			<=			16'h98B3;
		end
		32'h0000ED22: begin
				q			<=			16'h00D8;
		end
		32'h0000ED24: begin
				q			<=			16'hE5B3;
		end
		32'h0000ED26: begin
				q			<=			16'h0115;
		end
		32'h0000ED28: begin
				q			<=			16'hA823;
		end
		32'h0000ED2A: begin
				q			<=			16'h00B7;
		end
		32'h0000ED2C: begin
				q			<=			16'hF06F;
		end
		32'h0000ED2E: begin
				q			<=			16'hF4DF;
		end
		32'h0000ED30: begin
				q			<=			16'h87B7;
		end
		32'h0000ED32: begin
				q			<=			16'h0000;
		end
		32'h0000ED34: begin
				q			<=			16'h0863;
		end
		32'h0000ED36: begin
				q			<=			16'h0205;
		end
		32'h0000ED38: begin
				q			<=			16'h1793;
		end
		32'h0000ED3A: begin
				q			<=			16'h01C7;
		end
		32'h0000ED3C: begin
				q			<=			16'hD693;
		end
		32'h0000ED3E: begin
				q			<=			16'h0045;
		end
		32'h0000ED40: begin
				q			<=			16'hE7B3;
		end
		32'h0000ED42: begin
				q			<=			16'h00D7;
		end
		32'h0000ED44: begin
				q			<=			16'h2C23;
		end
		32'h0000ED46: begin
				q			<=			16'h00F1;
		end
		32'h0000ED48: begin
				q			<=			16'h5713;
		end
		32'h0000ED4A: begin
				q			<=			16'h0047;
		end
		32'h0000ED4C: begin
				q			<=			16'h87B7;
		end
		32'h0000ED4E: begin
				q			<=			16'h0000;
		end
		32'h0000ED50: begin
				q			<=			16'h9593;
		end
		32'h0000ED52: begin
				q			<=			16'h01C5;
		end
		32'h0000ED54: begin
				q			<=			16'h6733;
		end
		32'h0000ED56: begin
				q			<=			16'h00F7;
		end
		32'h0000ED58: begin
				q			<=			16'h2A23;
		end
		32'h0000ED5A: begin
				q			<=			16'h00B1;
		end
		32'h0000ED5C: begin
				q			<=			16'h2823;
		end
		32'h0000ED5E: begin
				q			<=			16'h0001;
		end
		32'h0000ED60: begin
				q			<=			16'h2E23;
		end
		32'h0000ED62: begin
				q			<=			16'h00E1;
		end
		32'h0000ED64: begin
				q			<=			16'h8793;
		end
		32'h0000ED66: begin
				q			<=			16'hFFF7;
		end
		32'h0000ED68: begin
				q			<=			16'hF06F;
		end
		32'h0000ED6A: begin
				q			<=			16'hE5DF;
		end
		32'h0000ED6C: begin
				q			<=			16'h0000;
		end
		32'h0000ED6E: begin
				q			<=			16'h0000;
		end
		32'h0000ED70: begin
				q			<=			16'h2583;
		end
		32'h0000ED72: begin
				q			<=			16'h00C5;
		end
		32'h0000ED74: begin
				q			<=			16'h2783;
		end
		32'h0000ED76: begin
				q			<=			16'h0085;
		end
		32'h0000ED78: begin
				q			<=			16'h2703;
		end
		32'h0000ED7A: begin
				q			<=			16'h0045;
		end
		32'h0000ED7C: begin
				q			<=			16'h0113;
		end
		32'h0000ED7E: begin
				q			<=			16'hFE01;
		end
		32'h0000ED80: begin
				q			<=			16'h2683;
		end
		32'h0000ED82: begin
				q			<=			16'h0005;
		end
		32'h0000ED84: begin
				q			<=			16'h2423;
		end
		32'h0000ED86: begin
				q			<=			16'h00F1;
		end
		32'h0000ED88: begin
				q			<=			16'h2C23;
		end
		32'h0000ED8A: begin
				q			<=			16'h00F1;
		end
		32'h0000ED8C: begin
				q			<=			16'h9793;
		end
		32'h0000ED8E: begin
				q			<=			16'h0105;
		end
		32'h0000ED90: begin
				q			<=			16'h2223;
		end
		32'h0000ED92: begin
				q			<=			16'h00E1;
		end
		32'h0000ED94: begin
				q			<=			16'h2A23;
		end
		32'h0000ED96: begin
				q			<=			16'h00E1;
		end
		32'h0000ED98: begin
				q			<=			16'hD793;
		end
		32'h0000ED9A: begin
				q			<=			16'h0107;
		end
		32'h0000ED9C: begin
				q			<=			16'h9713;
		end
		32'h0000ED9E: begin
				q			<=			16'h0015;
		end
		32'h0000EDA0: begin
				q			<=			16'h2623;
		end
		32'h0000EDA2: begin
				q			<=			16'h00B1;
		end
		32'h0000EDA4: begin
				q			<=			16'h2023;
		end
		32'h0000EDA6: begin
				q			<=			16'h00D1;
		end
		32'h0000EDA8: begin
				q			<=			16'h2823;
		end
		32'h0000EDAA: begin
				q			<=			16'h00D1;
		end
		32'h0000EDAC: begin
				q			<=			16'h2E23;
		end
		32'h0000EDAE: begin
				q			<=			16'h00F1;
		end
		32'h0000EDB0: begin
				q			<=			16'h5713;
		end
		32'h0000EDB2: begin
				q			<=			16'h0117;
		end
		32'h0000EDB4: begin
				q			<=			16'hD593;
		end
		32'h0000EDB6: begin
				q			<=			16'h01F5;
		end
		32'h0000EDB8: begin
				q			<=			16'h0313;
		end
		32'h0000EDBA: begin
				q			<=			16'h0101;
		end
		32'h0000EDBC: begin
				q			<=			16'h0613;
		end
		32'h0000EDBE: begin
				q			<=			16'h01C1;
		end
		32'h0000EDC0: begin
				q			<=			16'h2783;
		end
		32'h0000EDC2: begin
				q			<=			16'h0006;
		end
		32'h0000EDC4: begin
				q			<=			16'h2683;
		end
		32'h0000EDC6: begin
				q			<=			16'hFFC6;
		end
		32'h0000EDC8: begin
				q			<=			16'h0613;
		end
		32'h0000EDCA: begin
				q			<=			16'hFFC6;
		end
		32'h0000EDCC: begin
				q			<=			16'h9793;
		end
		32'h0000EDCE: begin
				q			<=			16'h0037;
		end
		32'h0000EDD0: begin
				q			<=			16'hD693;
		end
		32'h0000EDD2: begin
				q			<=			16'h01D6;
		end
		32'h0000EDD4: begin
				q			<=			16'hE7B3;
		end
		32'h0000EDD6: begin
				q			<=			16'h00D7;
		end
		32'h0000EDD8: begin
				q			<=			16'h2223;
		end
		32'h0000EDDA: begin
				q			<=			16'h00F6;
		end
		32'h0000EDDC: begin
				q			<=			16'h12E3;
		end
		32'h0000EDDE: begin
				q			<=			16'hFEC3;
		end
		32'h0000EDE0: begin
				q			<=			16'h2683;
		end
		32'h0000EDE2: begin
				q			<=			16'h0101;
		end
		32'h0000EDE4: begin
				q			<=			16'h0793;
		end
		32'h0000EDE6: begin
				q			<=			16'h0017;
		end
		32'h0000EDE8: begin
				q			<=			16'h9513;
		end
		32'h0000EDEA: begin
				q			<=			16'h0036;
		end
		32'h0000EDEC: begin
				q			<=			16'h86B7;
		end
		32'h0000EDEE: begin
				q			<=			16'h0000;
		end
		32'h0000EDF0: begin
				q			<=			16'h8693;
		end
		32'h0000EDF2: begin
				q			<=			16'hFFF6;
		end
		32'h0000EDF4: begin
				q			<=			16'hF7B3;
		end
		32'h0000EDF6: begin
				q			<=			16'h00D7;
		end
		32'h0000EDF8: begin
				q			<=			16'h2823;
		end
		32'h0000EDFA: begin
				q			<=			16'h00A1;
		end
		32'h0000EDFC: begin
				q			<=			16'h0693;
		end
		32'h0000EDFE: begin
				q			<=			16'h0010;
		end
		32'h0000EE00: begin
				q			<=			16'hDC63;
		end
		32'h0000EE02: begin
				q			<=			16'h1AF6;
		end
		32'h0000EE04: begin
				q			<=			16'hC7B7;
		end
		32'h0000EE06: begin
				q			<=			16'hFFFF;
		end
		32'h0000EE08: begin
				q			<=			16'h8793;
		end
		32'h0000EE0A: begin
				q			<=			16'h4007;
		end
		32'h0000EE0C: begin
				q			<=			16'h0733;
		end
		32'h0000EE0E: begin
				q			<=			16'h00F7;
		end
		32'h0000EE10: begin
				q			<=			16'h0793;
		end
		32'h0000EE12: begin
				q			<=			16'h7FE0;
		end
		32'h0000EE14: begin
				q			<=			16'hCE63;
		end
		32'h0000EE16: begin
				q			<=			16'h1EE7;
		end
		32'h0000EE18: begin
				q			<=			16'h5863;
		end
		32'h0000EE1A: begin
				q			<=			16'h06E0;
		end
		32'h0000EE1C: begin
				q			<=			16'h2783;
		end
		32'h0000EE1E: begin
				q			<=			16'h0181;
		end
		32'h0000EE20: begin
				q			<=			16'h2603;
		end
		32'h0000EE22: begin
				q			<=			16'h01C1;
		end
		32'h0000EE24: begin
				q			<=			16'h2803;
		end
		32'h0000EE26: begin
				q			<=			16'h0141;
		end
		32'h0000EE28: begin
				q			<=			16'hD693;
		end
		32'h0000EE2A: begin
				q			<=			16'h01C7;
		end
		32'h0000EE2C: begin
				q			<=			16'h1613;
		end
		32'h0000EE2E: begin
				q			<=			16'h0046;
		end
		32'h0000EE30: begin
				q			<=			16'h6633;
		end
		32'h0000EE32: begin
				q			<=			16'h00D6;
		end
		32'h0000EE34: begin
				q			<=			16'h1693;
		end
		32'h0000EE36: begin
				q			<=			16'h0048;
		end
		32'h0000EE38: begin
				q			<=			16'hE6B3;
		end
		32'h0000EE3A: begin
				q			<=			16'h00A6;
		end
		32'h0000EE3C: begin
				q			<=			16'h9793;
		end
		32'h0000EE3E: begin
				q			<=			16'h0047;
		end
		32'h0000EE40: begin
				q			<=			16'h5813;
		end
		32'h0000EE42: begin
				q			<=			16'h01C8;
		end
		32'h0000EE44: begin
				q			<=			16'h36B3;
		end
		32'h0000EE46: begin
				q			<=			16'h00D0;
		end
		32'h0000EE48: begin
				q			<=			16'hE7B3;
		end
		32'h0000EE4A: begin
				q			<=			16'h0107;
		end
		32'h0000EE4C: begin
				q			<=			16'hE6B3;
		end
		32'h0000EE4E: begin
				q			<=			16'h00F6;
		end
		32'h0000EE50: begin
				q			<=			16'h2A23;
		end
		32'h0000EE52: begin
				q			<=			16'h00C1;
		end
		32'h0000EE54: begin
				q			<=			16'h2823;
		end
		32'h0000EE56: begin
				q			<=			16'h00D1;
		end
		32'h0000EE58: begin
				q			<=			16'h2683;
		end
		32'h0000EE5A: begin
				q			<=			16'h0101;
		end
		32'h0000EE5C: begin
				q			<=			16'h2783;
		end
		32'h0000EE5E: begin
				q			<=			16'h0141;
		end
		32'h0000EE60: begin
				q			<=			16'hF613;
		end
		32'h0000EE62: begin
				q			<=			16'h0076;
		end
		32'h0000EE64: begin
				q			<=			16'h0C63;
		end
		32'h0000EE66: begin
				q			<=			16'h1A06;
		end
		32'h0000EE68: begin
				q			<=			16'hF613;
		end
		32'h0000EE6A: begin
				q			<=			16'h00F6;
		end
		32'h0000EE6C: begin
				q			<=			16'h0513;
		end
		32'h0000EE6E: begin
				q			<=			16'h0040;
		end
		32'h0000EE70: begin
				q			<=			16'h0663;
		end
		32'h0000EE72: begin
				q			<=			16'h1AA6;
		end
		32'h0000EE74: begin
				q			<=			16'h8613;
		end
		32'h0000EE76: begin
				q			<=			16'h0046;
		end
		32'h0000EE78: begin
				q			<=			16'h36B3;
		end
		32'h0000EE7A: begin
				q			<=			16'h00D6;
		end
		32'h0000EE7C: begin
				q			<=			16'h87B3;
		end
		32'h0000EE7E: begin
				q			<=			16'h00D7;
		end
		32'h0000EE80: begin
				q			<=			16'h0693;
		end
		32'h0000EE82: begin
				q			<=			16'h0006;
		end
		32'h0000EE84: begin
				q			<=			16'h006F;
		end
		32'h0000EE86: begin
				q			<=			16'h1980;
		end
		32'h0000EE88: begin
				q			<=			16'h0793;
		end
		32'h0000EE8A: begin
				q			<=			16'hFCC0;
		end
		32'h0000EE8C: begin
				q			<=			16'h5A63;
		end
		32'h0000EE8E: begin
				q			<=			16'h00F7;
		end
		32'h0000EE90: begin
				q			<=			16'h2A23;
		end
		32'h0000EE92: begin
				q			<=			16'h0001;
		end
		32'h0000EE94: begin
				q			<=			16'h2823;
		end
		32'h0000EE96: begin
				q			<=			16'h00D1;
		end
		32'h0000EE98: begin
				q			<=			16'h0713;
		end
		32'h0000EE9A: begin
				q			<=			16'h0000;
		end
		32'h0000EE9C: begin
				q			<=			16'hF06F;
		end
		32'h0000EE9E: begin
				q			<=			16'hFBDF;
		end
		32'h0000EEA0: begin
				q			<=			16'h2783;
		end
		32'h0000EEA2: begin
				q			<=			16'h01C1;
		end
		32'h0000EEA4: begin
				q			<=			16'h06B7;
		end
		32'h0000EEA6: begin
				q			<=			16'h0008;
		end
		32'h0000EEA8: begin
				q			<=			16'h0893;
		end
		32'h0000EEAA: begin
				q			<=			16'h0000;
		end
		32'h0000EEAC: begin
				q			<=			16'hE7B3;
		end
		32'h0000EEAE: begin
				q			<=			16'h00D7;
		end
		32'h0000EEB0: begin
				q			<=			16'h2E23;
		end
		32'h0000EEB2: begin
				q			<=			16'h00F1;
		end
		32'h0000EEB4: begin
				q			<=			16'h0793;
		end
		32'h0000EEB6: begin
				q			<=			16'h03D0;
		end
		32'h0000EEB8: begin
				q			<=			16'h8733;
		end
		32'h0000EEBA: begin
				q			<=			16'h40E7;
		end
		32'h0000EEBC: begin
				q			<=			16'h5513;
		end
		32'h0000EEBE: begin
				q			<=			16'h4057;
		end
		32'h0000EEC0: begin
				q			<=			16'h0793;
		end
		32'h0000EEC2: begin
				q			<=			16'h0003;
		end
		32'h0000EEC4: begin
				q			<=			16'h7713;
		end
		32'h0000EEC6: begin
				q			<=			16'h01F7;
		end
		32'h0000EEC8: begin
				q			<=			16'h0693;
		end
		32'h0000EECA: begin
				q			<=			16'h0000;
		end
		32'h0000EECC: begin
				q			<=			16'hA803;
		end
		32'h0000EECE: begin
				q			<=			16'h0007;
		end
		32'h0000EED0: begin
				q			<=			16'h8693;
		end
		32'h0000EED2: begin
				q			<=			16'h0016;
		end
		32'h0000EED4: begin
				q			<=			16'h8793;
		end
		32'h0000EED6: begin
				q			<=			16'h0047;
		end
		32'h0000EED8: begin
				q			<=			16'hE8B3;
		end
		32'h0000EEDA: begin
				q			<=			16'h0108;
		end
		32'h0000EEDC: begin
				q			<=			16'h18E3;
		end
		32'h0000EEDE: begin
				q			<=			16'hFED5;
		end
		32'h0000EEE0: begin
				q			<=			16'h9E93;
		end
		32'h0000EEE2: begin
				q			<=			16'h0026;
		end
		32'h0000EEE4: begin
				q			<=			16'h1E63;
		end
		32'h0000EEE6: begin
				q			<=			16'h0407;
		end
		32'h0000EEE8: begin
				q			<=			16'h0793;
		end
		32'h0000EEEA: begin
				q			<=			16'h0030;
		end
		32'h0000EEEC: begin
				q			<=			16'h87B3;
		end
		32'h0000EEEE: begin
				q			<=			16'h40D7;
		end
		32'h0000EEF0: begin
				q			<=			16'hDC63;
		end
		32'h0000EEF2: begin
				q			<=			16'h02E7;
		end
		32'h0000EEF4: begin
				q			<=			16'h0793;
		end
		32'h0000EEF6: begin
				q			<=			16'h0040;
		end
		32'h0000EEF8: begin
				q			<=			16'h86B3;
		end
		32'h0000EEFA: begin
				q			<=			16'h40D7;
		end
		32'h0000EEFC: begin
				q			<=			16'h0713;
		end
		32'h0000EEFE: begin
				q			<=			16'h0040;
		end
		32'h0000EF00: begin
				q			<=			16'h9793;
		end
		32'h0000EF02: begin
				q			<=			16'h0026;
		end
		32'h0000EF04: begin
				q			<=			16'h07B3;
		end
		32'h0000EF06: begin
				q			<=			16'h00F3;
		end
		32'h0000EF08: begin
				q			<=			16'hA023;
		end
		32'h0000EF0A: begin
				q			<=			16'h0007;
		end
		32'h0000EF0C: begin
				q			<=			16'h8693;
		end
		32'h0000EF0E: begin
				q			<=			16'h0016;
		end
		32'h0000EF10: begin
				q			<=			16'h98E3;
		end
		32'h0000EF12: begin
				q			<=			16'hFEE6;
		end
		32'h0000EF14: begin
				q			<=			16'h2703;
		end
		32'h0000EF16: begin
				q			<=			16'h0101;
		end
		32'h0000EF18: begin
				q			<=			16'h37B3;
		end
		32'h0000EF1A: begin
				q			<=			16'h0110;
		end
		32'h0000EF1C: begin
				q			<=			16'h67B3;
		end
		32'h0000EF1E: begin
				q			<=			16'h00F7;
		end
		32'h0000EF20: begin
				q			<=			16'h2823;
		end
		32'h0000EF22: begin
				q			<=			16'h00F1;
		end
		32'h0000EF24: begin
				q			<=			16'hF06F;
		end
		32'h0000EF26: begin
				q			<=			16'hF75F;
		end
		32'h0000EF28: begin
				q			<=			16'h0533;
		end
		32'h0000EF2A: begin
				q			<=			16'h01D6;
		end
		32'h0000EF2C: begin
				q			<=			16'h2503;
		end
		32'h0000EF2E: begin
				q			<=			16'h0005;
		end
		32'h0000EF30: begin
				q			<=			16'h0713;
		end
		32'h0000EF32: begin
				q			<=			16'h0017;
		end
		32'h0000EF34: begin
				q			<=			16'h0613;
		end
		32'h0000EF36: begin
				q			<=			16'h0046;
		end
		32'h0000EF38: begin
				q			<=			16'h2E23;
		end
		32'h0000EF3A: begin
				q			<=			16'hFEA6;
		end
		32'h0000EF3C: begin
				q			<=			16'hF06F;
		end
		32'h0000EF3E: begin
				q			<=			16'hFB5F;
		end
		32'h0000EF40: begin
				q			<=			16'h0793;
		end
		32'h0000EF42: begin
				q			<=			16'h0201;
		end
		32'h0000EF44: begin
				q			<=			16'h87B3;
		end
		32'h0000EF46: begin
				q			<=			16'h01D7;
		end
		32'h0000EF48: begin
				q			<=			16'hA783;
		end
		32'h0000EF4A: begin
				q			<=			16'hFF07;
		end
		32'h0000EF4C: begin
				q			<=			16'h0813;
		end
		32'h0000EF4E: begin
				q			<=			16'h0200;
		end
		32'h0000EF50: begin
				q			<=			16'h0833;
		end
		32'h0000EF52: begin
				q			<=			16'h40E8;
		end
		32'h0000EF54: begin
				q			<=			16'h97B3;
		end
		32'h0000EF56: begin
				q			<=			16'h0107;
		end
		32'h0000EF58: begin
				q			<=			16'hE8B3;
		end
		32'h0000EF5A: begin
				q			<=			16'h00F8;
		end
		32'h0000EF5C: begin
				q			<=			16'h0793;
		end
		32'h0000EF5E: begin
				q			<=			16'h0030;
		end
		32'h0000EF60: begin
				q			<=			16'h0E13;
		end
		32'h0000EF62: begin
				q			<=			16'h0000;
		end
		32'h0000EF64: begin
				q			<=			16'h87B3;
		end
		32'h0000EF66: begin
				q			<=			16'h40D7;
		end
		32'h0000EF68: begin
				q			<=			16'h4463;
		end
		32'h0000EF6A: begin
				q			<=			16'h02FE;
		end
		32'h0000EF6C: begin
				q			<=			16'h0613;
		end
		32'h0000EF6E: begin
				q			<=			16'h0040;
		end
		32'h0000EF70: begin
				q			<=			16'h06B3;
		end
		32'h0000EF72: begin
				q			<=			16'h40D6;
		end
		32'h0000EF74: begin
				q			<=			16'h9793;
		end
		32'h0000EF76: begin
				q			<=			16'h0027;
		end
		32'h0000EF78: begin
				q			<=			16'h0613;
		end
		32'h0000EF7A: begin
				q			<=			16'h0201;
		end
		32'h0000EF7C: begin
				q			<=			16'h07B3;
		end
		32'h0000EF7E: begin
				q			<=			16'h00F6;
		end
		32'h0000EF80: begin
				q			<=			16'h2603;
		end
		32'h0000EF82: begin
				q			<=			16'h01C1;
		end
		32'h0000EF84: begin
				q			<=			16'h5733;
		end
		32'h0000EF86: begin
				q			<=			16'h00E6;
		end
		32'h0000EF88: begin
				q			<=			16'hA823;
		end
		32'h0000EF8A: begin
				q			<=			16'hFEE7;
		end
		32'h0000EF8C: begin
				q			<=			16'hF06F;
		end
		32'h0000EF8E: begin
				q			<=			16'hF71F;
		end
		32'h0000EF90: begin
				q			<=			16'h0F33;
		end
		32'h0000EF92: begin
				q			<=			16'h01D6;
		end
		32'h0000EF94: begin
				q			<=			16'h2503;
		end
		32'h0000EF96: begin
				q			<=			16'h000F;
		end
		32'h0000EF98: begin
				q			<=			16'h2F03;
		end
		32'h0000EF9A: begin
				q			<=			16'h004F;
		end
		32'h0000EF9C: begin
				q			<=			16'h0E13;
		end
		32'h0000EF9E: begin
				q			<=			16'h001E;
		end
		32'h0000EFA0: begin
				q			<=			16'h5533;
		end
		32'h0000EFA2: begin
				q			<=			16'h00E5;
		end
		32'h0000EFA4: begin
				q			<=			16'h1F33;
		end
		32'h0000EFA6: begin
				q			<=			16'h010F;
		end
		32'h0000EFA8: begin
				q			<=			16'h6533;
		end
		32'h0000EFAA: begin
				q			<=			16'h01E5;
		end
		32'h0000EFAC: begin
				q			<=			16'h2023;
		end
		32'h0000EFAE: begin
				q			<=			16'h00A6;
		end
		32'h0000EFB0: begin
				q			<=			16'h0613;
		end
		32'h0000EFB2: begin
				q			<=			16'h0046;
		end
		32'h0000EFB4: begin
				q			<=			16'hF06F;
		end
		32'h0000EFB6: begin
				q			<=			16'hFB5F;
		end
		32'h0000EFB8: begin
				q			<=			16'h2603;
		end
		32'h0000EFBA: begin
				q			<=			16'h0141;
		end
		32'h0000EFBC: begin
				q			<=			16'h2783;
		end
		32'h0000EFBE: begin
				q			<=			16'h0181;
		end
		32'h0000EFC0: begin
				q			<=			16'h2803;
		end
		32'h0000EFC2: begin
				q			<=			16'h01C1;
		end
		32'h0000EFC4: begin
				q			<=			16'h66B3;
		end
		32'h0000EFC6: begin
				q			<=			16'h00F6;
		end
		32'h0000EFC8: begin
				q			<=			16'hE6B3;
		end
		32'h0000EFCA: begin
				q			<=			16'h0106;
		end
		32'h0000EFCC: begin
				q			<=			16'hE6B3;
		end
		32'h0000EFCE: begin
				q			<=			16'h00A6;
		end
		32'h0000EFD0: begin
				q			<=			16'h1863;
		end
		32'h0000EFD2: begin
				q			<=			16'h0007;
		end
		32'h0000EFD4: begin
				q			<=			16'h36B3;
		end
		32'h0000EFD6: begin
				q			<=			16'h00D0;
		end
		32'h0000EFD8: begin
				q			<=			16'h0793;
		end
		32'h0000EFDA: begin
				q			<=			16'h0000;
		end
		32'h0000EFDC: begin
				q			<=			16'hF06F;
		end
		32'h0000EFDE: begin
				q			<=			16'hE85F;
		end
		32'h0000EFE0: begin
				q			<=			16'h8A63;
		end
		32'h0000EFE2: begin
				q			<=			16'h0C06;
		end
		32'h0000EFE4: begin
				q			<=			16'h5693;
		end
		32'h0000EFE6: begin
				q			<=			16'h01C6;
		end
		32'h0000EFE8: begin
				q			<=			16'h1813;
		end
		32'h0000EFEA: begin
				q			<=			16'h0048;
		end
		32'h0000EFEC: begin
				q			<=			16'h9613;
		end
		32'h0000EFEE: begin
				q			<=			16'h0047;
		end
		32'h0000EFF0: begin
				q			<=			16'hD793;
		end
		32'h0000EFF2: begin
				q			<=			16'h01C7;
		end
		32'h0000EFF4: begin
				q			<=			16'h0737;
		end
		32'h0000EFF6: begin
				q			<=			16'h0040;
		end
		32'h0000EFF8: begin
				q			<=			16'hE6B3;
		end
		32'h0000EFFA: begin
				q			<=			16'h00C6;
		end
		32'h0000EFFC: begin
				q			<=			16'hE7B3;
		end
		32'h0000EFFE: begin
				q			<=			16'h0107;
		end
		32'h0000F000: begin
				q			<=			16'hE7B3;
		end
		32'h0000F002: begin
				q			<=			16'h00E7;
		end
		32'h0000F004: begin
				q			<=			16'hF693;
		end
		32'h0000F006: begin
				q			<=			16'hFF86;
		end
		32'h0000F008: begin
				q			<=			16'h0713;
		end
		32'h0000F00A: begin
				q			<=			16'h7FF0;
		end
		32'h0000F00C: begin
				q			<=			16'hF06F;
		end
		32'h0000F00E: begin
				q			<=			16'hE55F;
		end
		32'h0000F010: begin
				q			<=			16'h0793;
		end
		32'h0000F012: begin
				q			<=			16'h0000;
		end
		32'h0000F014: begin
				q			<=			16'h0693;
		end
		32'h0000F016: begin
				q			<=			16'h0000;
		end
		32'h0000F018: begin
				q			<=			16'h0713;
		end
		32'h0000F01A: begin
				q			<=			16'h7FF0;
		end
		32'h0000F01C: begin
				q			<=			16'h9613;
		end
		32'h0000F01E: begin
				q			<=			16'h0087;
		end
		32'h0000F020: begin
				q			<=			16'h5E63;
		end
		32'h0000F022: begin
				q			<=			16'h0006;
		end
		32'h0000F024: begin
				q			<=			16'h0713;
		end
		32'h0000F026: begin
				q			<=			16'h0017;
		end
		32'h0000F028: begin
				q			<=			16'h0613;
		end
		32'h0000F02A: begin
				q			<=			16'h7FF0;
		end
		32'h0000F02C: begin
				q			<=			16'h0863;
		end
		32'h0000F02E: begin
				q			<=			16'h08C7;
		end
		32'h0000F030: begin
				q			<=			16'h0637;
		end
		32'h0000F032: begin
				q			<=			16'hFF80;
		end
		32'h0000F034: begin
				q			<=			16'h0613;
		end
		32'h0000F036: begin
				q			<=			16'hFFF6;
		end
		32'h0000F038: begin
				q			<=			16'hF7B3;
		end
		32'h0000F03A: begin
				q			<=			16'h00C7;
		end
		32'h0000F03C: begin
				q			<=			16'h9613;
		end
		32'h0000F03E: begin
				q			<=			16'h01D7;
		end
		32'h0000F040: begin
				q			<=			16'hD693;
		end
		32'h0000F042: begin
				q			<=			16'h0036;
		end
		32'h0000F044: begin
				q			<=			16'h66B3;
		end
		32'h0000F046: begin
				q			<=			16'h00D6;
		end
		32'h0000F048: begin
				q			<=			16'h0613;
		end
		32'h0000F04A: begin
				q			<=			16'h7FF0;
		end
		32'h0000F04C: begin
				q			<=			16'hD793;
		end
		32'h0000F04E: begin
				q			<=			16'h0037;
		end
		32'h0000F050: begin
				q			<=			16'h1E63;
		end
		32'h0000F052: begin
				q			<=			16'h00C7;
		end
		32'h0000F054: begin
				q			<=			16'hE6B3;
		end
		32'h0000F056: begin
				q			<=			16'h00F6;
		end
		32'h0000F058: begin
				q			<=			16'h0793;
		end
		32'h0000F05A: begin
				q			<=			16'h0000;
		end
		32'h0000F05C: begin
				q			<=			16'h8863;
		end
		32'h0000F05E: begin
				q			<=			16'h0006;
		end
		32'h0000F060: begin
				q			<=			16'h07B7;
		end
		32'h0000F062: begin
				q			<=			16'h0008;
		end
		32'h0000F064: begin
				q			<=			16'h0693;
		end
		32'h0000F066: begin
				q			<=			16'h0000;
		end
		32'h0000F068: begin
				q			<=			16'h0593;
		end
		32'h0000F06A: begin
				q			<=			16'h0000;
		end
		32'h0000F06C: begin
				q			<=			16'h0637;
		end
		32'h0000F06E: begin
				q			<=			16'h0010;
		end
		32'h0000F070: begin
				q			<=			16'h0613;
		end
		32'h0000F072: begin
				q			<=			16'hFFF6;
		end
		32'h0000F074: begin
				q			<=			16'hF7B3;
		end
		32'h0000F076: begin
				q			<=			16'h00C7;
		end
		32'h0000F078: begin
				q			<=			16'h0637;
		end
		32'h0000F07A: begin
				q			<=			16'h8010;
		end
		32'h0000F07C: begin
				q			<=			16'h7713;
		end
		32'h0000F07E: begin
				q			<=			16'h7FF7;
		end
		32'h0000F080: begin
				q			<=			16'h0613;
		end
		32'h0000F082: begin
				q			<=			16'hFFF6;
		end
		32'h0000F084: begin
				q			<=			16'h1713;
		end
		32'h0000F086: begin
				q			<=			16'h0147;
		end
		32'h0000F088: begin
				q			<=			16'hF7B3;
		end
		32'h0000F08A: begin
				q			<=			16'h00C7;
		end
		32'h0000F08C: begin
				q			<=			16'hE7B3;
		end
		32'h0000F08E: begin
				q			<=			16'h00E7;
		end
		32'h0000F090: begin
				q			<=			16'h0737;
		end
		32'h0000F092: begin
				q			<=			16'h8000;
		end
		32'h0000F094: begin
				q			<=			16'h4713;
		end
		32'h0000F096: begin
				q			<=			16'hFFF7;
		end
		32'h0000F098: begin
				q			<=			16'h9593;
		end
		32'h0000F09A: begin
				q			<=			16'h01F5;
		end
		32'h0000F09C: begin
				q			<=			16'hF7B3;
		end
		32'h0000F09E: begin
				q			<=			16'h00E7;
		end
		32'h0000F0A0: begin
				q			<=			16'hE733;
		end
		32'h0000F0A2: begin
				q			<=			16'h00B7;
		end
		32'h0000F0A4: begin
				q			<=			16'h8513;
		end
		32'h0000F0A6: begin
				q			<=			16'h0006;
		end
		32'h0000F0A8: begin
				q			<=			16'h0593;
		end
		32'h0000F0AA: begin
				q			<=			16'h0007;
		end
		32'h0000F0AC: begin
				q			<=			16'h0113;
		end
		32'h0000F0AE: begin
				q			<=			16'h0201;
		end
		32'h0000F0B0: begin
				q			<=			16'h8067;
		end
		32'h0000F0B2: begin
				q			<=			16'h0000;
		end
		32'h0000F0B4: begin
				q			<=			16'h0793;
		end
		32'h0000F0B6: begin
				q			<=			16'h0000;
		end
		32'h0000F0B8: begin
				q			<=			16'hF06F;
		end
		32'h0000F0BA: begin
				q			<=			16'hF61F;
		end
		32'h0000F0BC: begin
				q			<=			16'h0793;
		end
		32'h0000F0BE: begin
				q			<=			16'h0000;
		end
		32'h0000F0C0: begin
				q			<=			16'h0693;
		end
		32'h0000F0C2: begin
				q			<=			16'h0000;
		end
		32'h0000F0C4: begin
				q			<=			16'hF06F;
		end
		32'h0000F0C6: begin
				q			<=			16'hF79F;
		end
		32'h0000F0C8: begin
				q			<=			16'h0000;
		end
		32'h0000F0CA: begin
				q			<=			16'h0000;
		end
		32'h0000F0CC: begin
				q			<=			16'h07B7;
		end
		32'h0000F0CE: begin
				q			<=			16'h0001;
		end
		32'h0000F0D0: begin
				q			<=			16'h7A63;
		end
		32'h0000F0D2: begin
				q			<=			16'h02F5;
		end
		32'h0000F0D4: begin
				q			<=			16'h0793;
		end
		32'h0000F0D6: begin
				q			<=			16'h0FF0;
		end
		32'h0000F0D8: begin
				q			<=			16'hB7B3;
		end
		32'h0000F0DA: begin
				q			<=			16'h00A7;
		end
		32'h0000F0DC: begin
				q			<=			16'h9793;
		end
		32'h0000F0DE: begin
				q			<=			16'h0037;
		end
		32'h0000F0E0: begin
				q			<=			16'h0713;
		end
		32'h0000F0E2: begin
				q			<=			16'h0200;
		end
		32'h0000F0E4: begin
				q			<=			16'h0733;
		end
		32'h0000F0E6: begin
				q			<=			16'h40F7;
		end
		32'h0000F0E8: begin
				q			<=			16'h57B3;
		end
		32'h0000F0EA: begin
				q			<=			16'h00F5;
		end
		32'h0000F0EC: begin
				q			<=			16'h1517;
		end
		32'h0000F0EE: begin
				q			<=			16'h0000;
		end
		32'h0000F0F0: begin
				q			<=			16'h0513;
		end
		32'h0000F0F2: begin
				q			<=			16'h8805;
		end
		32'h0000F0F4: begin
				q			<=			16'h07B3;
		end
		32'h0000F0F6: begin
				q			<=			16'h00F5;
		end
		32'h0000F0F8: begin
				q			<=			16'hC503;
		end
		32'h0000F0FA: begin
				q			<=			16'h0007;
		end
		32'h0000F0FC: begin
				q			<=			16'h0533;
		end
		32'h0000F0FE: begin
				q			<=			16'h40A7;
		end
		32'h0000F100: begin
				q			<=			16'h8067;
		end
		32'h0000F102: begin
				q			<=			16'h0000;
		end
		32'h0000F104: begin
				q			<=			16'h0737;
		end
		32'h0000F106: begin
				q			<=			16'h0100;
		end
		32'h0000F108: begin
				q			<=			16'h0793;
		end
		32'h0000F10A: begin
				q			<=			16'h0100;
		end
		32'h0000F10C: begin
				q			<=			16'h6AE3;
		end
		32'h0000F10E: begin
				q			<=			16'hFCE5;
		end
		32'h0000F110: begin
				q			<=			16'h0793;
		end
		32'h0000F112: begin
				q			<=			16'h0180;
		end
		32'h0000F114: begin
				q			<=			16'hF06F;
		end
		32'h0000F116: begin
				q			<=			16'hFCDF;
		end
		32'h0000F118: begin
				q			<=			16'h0000;
		end
		32'h0000F11A: begin
				q			<=			16'h0000;
		end
		32'h0000F11C: begin
				q			<=			16'h0000;
		end
		32'h0000F11E: begin
				q			<=			16'h0000;
		end
		32'h0000F120: begin
				q			<=			16'h4034;
		end
		32'h0000F122: begin
				q			<=			16'hFFFF;
		end
		32'h0000F124: begin
				q			<=			16'h51F8;
		end
		32'h0000F126: begin
				q			<=			16'hFFFF;
		end
		32'h0000F128: begin
				q			<=			16'h51F8;
		end
		32'h0000F12A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F12C: begin
				q			<=			16'h4048;
		end
		32'h0000F12E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F130: begin
				q			<=			16'h51F8;
		end
		32'h0000F132: begin
				q			<=			16'hFFFF;
		end
		32'h0000F134: begin
				q			<=			16'h51F8;
		end
		32'h0000F136: begin
				q			<=			16'hFFFF;
		end
		32'h0000F138: begin
				q			<=			16'h51F8;
		end
		32'h0000F13A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F13C: begin
				q			<=			16'h3FD8;
		end
		32'h0000F13E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F140: begin
				q			<=			16'h51F8;
		end
		32'h0000F142: begin
				q			<=			16'hFFFF;
		end
		32'h0000F144: begin
				q			<=			16'h51F8;
		end
		32'h0000F146: begin
				q			<=			16'hFFFF;
		end
		32'h0000F148: begin
				q			<=			16'h4050;
		end
		32'h0000F14A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F14C: begin
				q			<=			16'h4070;
		end
		32'h0000F14E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F150: begin
				q			<=			16'h51F8;
		end
		32'h0000F152: begin
				q			<=			16'hFFFF;
		end
		32'h0000F154: begin
				q			<=			16'h4068;
		end
		32'h0000F156: begin
				q			<=			16'hFFFF;
		end
		32'h0000F158: begin
				q			<=			16'h4078;
		end
		32'h0000F15A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F15C: begin
				q			<=			16'h51F8;
		end
		32'h0000F15E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F160: begin
				q			<=			16'h40D0;
		end
		32'h0000F162: begin
				q			<=			16'hFFFF;
		end
		32'h0000F164: begin
				q			<=			16'h40D8;
		end
		32'h0000F166: begin
				q			<=			16'hFFFF;
		end
		32'h0000F168: begin
				q			<=			16'h40D8;
		end
		32'h0000F16A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F16C: begin
				q			<=			16'h40D8;
		end
		32'h0000F16E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F170: begin
				q			<=			16'h40D8;
		end
		32'h0000F172: begin
				q			<=			16'hFFFF;
		end
		32'h0000F174: begin
				q			<=			16'h40D8;
		end
		32'h0000F176: begin
				q			<=			16'hFFFF;
		end
		32'h0000F178: begin
				q			<=			16'h40D8;
		end
		32'h0000F17A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F17C: begin
				q			<=			16'h40D8;
		end
		32'h0000F17E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F180: begin
				q			<=			16'h40D8;
		end
		32'h0000F182: begin
				q			<=			16'hFFFF;
		end
		32'h0000F184: begin
				q			<=			16'h40D8;
		end
		32'h0000F186: begin
				q			<=			16'hFFFF;
		end
		32'h0000F188: begin
				q			<=			16'h51F8;
		end
		32'h0000F18A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F18C: begin
				q			<=			16'h51F8;
		end
		32'h0000F18E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F190: begin
				q			<=			16'h51F8;
		end
		32'h0000F192: begin
				q			<=			16'hFFFF;
		end
		32'h0000F194: begin
				q			<=			16'h51F8;
		end
		32'h0000F196: begin
				q			<=			16'hFFFF;
		end
		32'h0000F198: begin
				q			<=			16'h51F8;
		end
		32'h0000F19A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F19C: begin
				q			<=			16'h51F8;
		end
		32'h0000F19E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1A0: begin
				q			<=			16'h51F8;
		end
		32'h0000F1A2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1A4: begin
				q			<=			16'h424C;
		end
		32'h0000F1A6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1A8: begin
				q			<=			16'h51F8;
		end
		32'h0000F1AA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1AC: begin
				q			<=			16'h416C;
		end
		32'h0000F1AE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1B0: begin
				q			<=			16'h41A0;
		end
		32'h0000F1B2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1B4: begin
				q			<=			16'h424C;
		end
		32'h0000F1B6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1B8: begin
				q			<=			16'h424C;
		end
		32'h0000F1BA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1BC: begin
				q			<=			16'h424C;
		end
		32'h0000F1BE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1C0: begin
				q			<=			16'h51F8;
		end
		32'h0000F1C2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1C4: begin
				q			<=			16'h51F8;
		end
		32'h0000F1C6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1C8: begin
				q			<=			16'h51F8;
		end
		32'h0000F1CA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1CC: begin
				q			<=			16'h51F8;
		end
		32'h0000F1CE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1D0: begin
				q			<=			16'h410C;
		end
		32'h0000F1D2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1D4: begin
				q			<=			16'h51F8;
		end
		32'h0000F1D6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1D8: begin
				q			<=			16'h51F8;
		end
		32'h0000F1DA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1DC: begin
				q			<=			16'h4BF0;
		end
		32'h0000F1DE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1E0: begin
				q			<=			16'h51F8;
		end
		32'h0000F1E2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1E4: begin
				q			<=			16'h51F8;
		end
		32'h0000F1E6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1E8: begin
				q			<=			16'h51F8;
		end
		32'h0000F1EA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1EC: begin
				q			<=			16'h4CBC;
		end
		32'h0000F1EE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1F0: begin
				q			<=			16'h51F8;
		end
		32'h0000F1F2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1F4: begin
				q			<=			16'h4FA0;
		end
		32'h0000F1F6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1F8: begin
				q			<=			16'h51F8;
		end
		32'h0000F1FA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F1FC: begin
				q			<=			16'h51F8;
		end
		32'h0000F1FE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F200: begin
				q			<=			16'h3F7C;
		end
		32'h0000F202: begin
				q			<=			16'hFFFF;
		end
		32'h0000F204: begin
				q			<=			16'h51F8;
		end
		32'h0000F206: begin
				q			<=			16'hFFFF;
		end
		32'h0000F208: begin
				q			<=			16'h51F8;
		end
		32'h0000F20A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F20C: begin
				q			<=			16'h51F8;
		end
		32'h0000F20E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F210: begin
				q			<=			16'h51F8;
		end
		32'h0000F212: begin
				q			<=			16'hFFFF;
		end
		32'h0000F214: begin
				q			<=			16'h51F8;
		end
		32'h0000F216: begin
				q			<=			16'hFFFF;
		end
		32'h0000F218: begin
				q			<=			16'h51F8;
		end
		32'h0000F21A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F21C: begin
				q			<=			16'h51F8;
		end
		32'h0000F21E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F220: begin
				q			<=			16'h51F8;
		end
		32'h0000F222: begin
				q			<=			16'hFFFF;
		end
		32'h0000F224: begin
				q			<=			16'h424C;
		end
		32'h0000F226: begin
				q			<=			16'hFFFF;
		end
		32'h0000F228: begin
				q			<=			16'h51F8;
		end
		32'h0000F22A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F22C: begin
				q			<=			16'h416C;
		end
		32'h0000F22E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F230: begin
				q			<=			16'h41A4;
		end
		32'h0000F232: begin
				q			<=			16'hFFFF;
		end
		32'h0000F234: begin
				q			<=			16'h424C;
		end
		32'h0000F236: begin
				q			<=			16'hFFFF;
		end
		32'h0000F238: begin
				q			<=			16'h424C;
		end
		32'h0000F23A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F23C: begin
				q			<=			16'h424C;
		end
		32'h0000F23E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F240: begin
				q			<=			16'h4114;
		end
		32'h0000F242: begin
				q			<=			16'hFFFF;
		end
		32'h0000F244: begin
				q			<=			16'h41A4;
		end
		32'h0000F246: begin
				q			<=			16'hFFFF;
		end
		32'h0000F248: begin
				q			<=			16'h415C;
		end
		32'h0000F24A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F24C: begin
				q			<=			16'h51F8;
		end
		32'h0000F24E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F250: begin
				q			<=			16'h4140;
		end
		32'h0000F252: begin
				q			<=			16'hFFFF;
		end
		32'h0000F254: begin
				q			<=			16'h51F8;
		end
		32'h0000F256: begin
				q			<=			16'hFFFF;
		end
		32'h0000F258: begin
				q			<=			16'h4B84;
		end
		32'h0000F25A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F25C: begin
				q			<=			16'h4BF4;
		end
		32'h0000F25E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F260: begin
				q			<=			16'h4C84;
		end
		32'h0000F262: begin
				q			<=			16'hFFFF;
		end
		32'h0000F264: begin
				q			<=			16'h415C;
		end
		32'h0000F266: begin
				q			<=			16'hFFFF;
		end
		32'h0000F268: begin
				q			<=			16'h51F8;
		end
		32'h0000F26A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F26C: begin
				q			<=			16'h4CBC;
		end
		32'h0000F26E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F270: begin
				q			<=			16'h3F3C;
		end
		32'h0000F272: begin
				q			<=			16'hFFFF;
		end
		32'h0000F274: begin
				q			<=			16'h4FA4;
		end
		32'h0000F276: begin
				q			<=			16'hFFFF;
		end
		32'h0000F278: begin
				q			<=			16'h51F8;
		end
		32'h0000F27A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F27C: begin
				q			<=			16'h51F8;
		end
		32'h0000F27E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F280: begin
				q			<=			16'h5008;
		end
		32'h0000F282: begin
				q			<=			16'hFFFF;
		end
		32'h0000F284: begin
				q			<=			16'h51F8;
		end
		32'h0000F286: begin
				q			<=			16'hFFFF;
		end
		32'h0000F288: begin
				q			<=			16'h3F3C;
		end
		32'h0000F28A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F28C: begin
				q			<=			16'h2020;
		end
		32'h0000F28E: begin
				q			<=			16'h2020;
		end
		32'h0000F290: begin
				q			<=			16'h2020;
		end
		32'h0000F292: begin
				q			<=			16'h2020;
		end
		32'h0000F294: begin
				q			<=			16'h2020;
		end
		32'h0000F296: begin
				q			<=			16'h2020;
		end
		32'h0000F298: begin
				q			<=			16'h2020;
		end
		32'h0000F29A: begin
				q			<=			16'h2020;
		end
		32'h0000F29C: begin
				q			<=			16'h3030;
		end
		32'h0000F29E: begin
				q			<=			16'h3030;
		end
		32'h0000F2A0: begin
				q			<=			16'h3030;
		end
		32'h0000F2A2: begin
				q			<=			16'h3030;
		end
		32'h0000F2A4: begin
				q			<=			16'h3030;
		end
		32'h0000F2A6: begin
				q			<=			16'h3030;
		end
		32'h0000F2A8: begin
				q			<=			16'h3030;
		end
		32'h0000F2AA: begin
				q			<=			16'h3030;
		end
		32'h0000F2AC: begin
				q			<=			16'h0000;
		end
		32'h0000F2AE: begin
				q			<=			16'h0000;
		end
		32'h0000F2B0: begin
				q			<=			16'h0000;
		end
		32'h0000F2B2: begin
				q			<=			16'h0000;
		end
		32'h0000F2B4: begin
				q			<=			16'h0000;
		end
		32'h0000F2B6: begin
				q			<=			16'h0000;
		end
		32'h0000F2B8: begin
				q			<=			16'h0000;
		end
		32'h0000F2BA: begin
				q			<=			16'h0000;
		end
		32'h0000F2BC: begin
				q			<=			16'h0000;
		end
		32'h0000F2BE: begin
				q			<=			16'h0000;
		end
		32'h0000F2C0: begin
				q			<=			16'h0000;
		end
		32'h0000F2C2: begin
				q			<=			16'h0000;
		end
		32'h0000F2C4: begin
				q			<=			16'h0000;
		end
		32'h0000F2C6: begin
				q			<=			16'h0000;
		end
		32'h0000F2C8: begin
				q			<=			16'h0000;
		end
		32'h0000F2CA: begin
				q			<=			16'h0000;
		end
		32'h0000F2CC: begin
				q			<=			16'h0000;
		end
		32'h0000F2CE: begin
				q			<=			16'h0000;
		end
		32'h0000F2D0: begin
				q			<=			16'h8000;
		end
		32'h0000F2D2: begin
				q			<=			16'h3FFF;
		end
		32'h0000F2D4: begin
				q			<=			16'h6576;
		end
		32'h0000F2D6: begin
				q			<=			16'h4A92;
		end
		32'h0000F2D8: begin
				q			<=			16'h804A;
		end
		32'h0000F2DA: begin
				q			<=			16'h153F;
		end
		32'h0000F2DC: begin
				q			<=			16'hC94C;
		end
		32'h0000F2DE: begin
				q			<=			16'h979A;
		end
		32'h0000F2E0: begin
				q			<=			16'h8A20;
		end
		32'h0000F2E2: begin
				q			<=			16'h5202;
		end
		32'h0000F2E4: begin
				q			<=			16'hC460;
		end
		32'h0000F2E6: begin
				q			<=			16'h7525;
		end
		32'h0000F2E8: begin
				q			<=			16'h6A32;
		end
		32'h0000F2EA: begin
				q			<=			16'hCE52;
		end
		32'h0000F2EC: begin
				q			<=			16'h329A;
		end
		32'h0000F2EE: begin
				q			<=			16'h28CE;
		end
		32'h0000F2F0: begin
				q			<=			16'hA74D;
		end
		32'h0000F2F2: begin
				q			<=			16'h5DE4;
		end
		32'h0000F2F4: begin
				q			<=			16'hC53D;
		end
		32'h0000F2F6: begin
				q			<=			16'h3B5D;
		end
		32'h0000F2F8: begin
				q			<=			16'h9E8B;
		end
		32'h0000F2FA: begin
				q			<=			16'h5A92;
		end
		32'h0000F2FC: begin
				q			<=			16'h526C;
		end
		32'h0000F2FE: begin
				q			<=			16'h50CE;
		end
		32'h0000F300: begin
				q			<=			16'hF18B;
		end
		32'h0000F302: begin
				q			<=			16'h3D28;
		end
		32'h0000F304: begin
				q			<=			16'h650D;
		end
		32'h0000F306: begin
				q			<=			16'h0C17;
		end
		32'h0000F308: begin
				q			<=			16'h8175;
		end
		32'h0000F30A: begin
				q			<=			16'h7586;
		end
		32'h0000F30C: begin
				q			<=			16'hC976;
		end
		32'h0000F30E: begin
				q			<=			16'h4D48;
		end
		32'h0000F310: begin
				q			<=			16'h9C66;
		end
		32'h0000F312: begin
				q			<=			16'h58F8;
		end
		32'h0000F314: begin
				q			<=			16'hBC50;
		end
		32'h0000F316: begin
				q			<=			16'h5C54;
		end
		32'h0000F318: begin
				q			<=			16'hCC65;
		end
		32'h0000F31A: begin
				q			<=			16'h91C6;
		end
		32'h0000F31C: begin
				q			<=			16'hA60E;
		end
		32'h0000F31E: begin
				q			<=			16'hA0AE;
		end
		32'h0000F320: begin
				q			<=			16'hE319;
		end
		32'h0000F322: begin
				q			<=			16'h46A3;
		end
		32'h0000F324: begin
				q			<=			16'h851E;
		end
		32'h0000F326: begin
				q			<=			16'hEAB7;
		end
		32'h0000F328: begin
				q			<=			16'h98FE;
		end
		32'h0000F32A: begin
				q			<=			16'h901B;
		end
		32'h0000F32C: begin
				q			<=			16'hDDBB;
		end
		32'h0000F32E: begin
				q			<=			16'hDE8D;
		end
		32'h0000F330: begin
				q			<=			16'h9DF9;
		end
		32'h0000F332: begin
				q			<=			16'hEBFB;
		end
		32'h0000F334: begin
				q			<=			16'hAA7E;
		end
		32'h0000F336: begin
				q			<=			16'h4351;
		end
		32'h0000F338: begin
				q			<=			16'h0235;
		end
		32'h0000F33A: begin
				q			<=			16'h0137;
		end
		32'h0000F33C: begin
				q			<=			16'h36B1;
		end
		32'h0000F33E: begin
				q			<=			16'h336C;
		end
		32'h0000F340: begin
				q			<=			16'hC66F;
		end
		32'h0000F342: begin
				q			<=			16'h8CDF;
		end
		32'h0000F344: begin
				q			<=			16'h80E9;
		end
		32'h0000F346: begin
				q			<=			16'h47C9;
		end
		32'h0000F348: begin
				q			<=			16'h93BA;
		end
		32'h0000F34A: begin
				q			<=			16'h41A8;
		end
		32'h0000F34C: begin
				q			<=			16'h50F8;
		end
		32'h0000F34E: begin
				q			<=			16'h25FB;
		end
		32'h0000F350: begin
				q			<=			16'hC76B;
		end
		32'h0000F352: begin
				q			<=			16'h6B71;
		end
		32'h0000F354: begin
				q			<=			16'h3CBF;
		end
		32'h0000F356: begin
				q			<=			16'hA6D5;
		end
		32'h0000F358: begin
				q			<=			16'hFFCF;
		end
		32'h0000F35A: begin
				q			<=			16'h1F49;
		end
		32'h0000F35C: begin
				q			<=			16'hC278;
		end
		32'h0000F35E: begin
				q			<=			16'h40D3;
		end
		32'h0000F360: begin
				q			<=			16'h0000;
		end
		32'h0000F362: begin
				q			<=			16'h0000;
		end
		32'h0000F364: begin
				q			<=			16'h0000;
		end
		32'h0000F366: begin
				q			<=			16'h0000;
		end
		32'h0000F368: begin
				q			<=			16'hF020;
		end
		32'h0000F36A: begin
				q			<=			16'hB59D;
		end
		32'h0000F36C: begin
				q			<=			16'h2B70;
		end
		32'h0000F36E: begin
				q			<=			16'hADA8;
		end
		32'h0000F370: begin
				q			<=			16'h9DC5;
		end
		32'h0000F372: begin
				q			<=			16'h4069;
		end
		32'h0000F374: begin
				q			<=			16'h0000;
		end
		32'h0000F376: begin
				q			<=			16'h0000;
		end
		32'h0000F378: begin
				q			<=			16'h0000;
		end
		32'h0000F37A: begin
				q			<=			16'h0000;
		end
		32'h0000F37C: begin
				q			<=			16'h0000;
		end
		32'h0000F37E: begin
				q			<=			16'h0000;
		end
		32'h0000F380: begin
				q			<=			16'h0400;
		end
		32'h0000F382: begin
				q			<=			16'hC9BF;
		end
		32'h0000F384: begin
				q			<=			16'h8E1B;
		end
		32'h0000F386: begin
				q			<=			16'h4034;
		end
		32'h0000F388: begin
				q			<=			16'h0000;
		end
		32'h0000F38A: begin
				q			<=			16'h0000;
		end
		32'h0000F38C: begin
				q			<=			16'h0000;
		end
		32'h0000F38E: begin
				q			<=			16'h0000;
		end
		32'h0000F390: begin
				q			<=			16'h0000;
		end
		32'h0000F392: begin
				q			<=			16'h0000;
		end
		32'h0000F394: begin
				q			<=			16'h0000;
		end
		32'h0000F396: begin
				q			<=			16'h2000;
		end
		32'h0000F398: begin
				q			<=			16'hBEBC;
		end
		32'h0000F39A: begin
				q			<=			16'h4019;
		end
		32'h0000F39C: begin
				q			<=			16'h0000;
		end
		32'h0000F39E: begin
				q			<=			16'h0000;
		end
		32'h0000F3A0: begin
				q			<=			16'h0000;
		end
		32'h0000F3A2: begin
				q			<=			16'h0000;
		end
		32'h0000F3A4: begin
				q			<=			16'h0000;
		end
		32'h0000F3A6: begin
				q			<=			16'h0000;
		end
		32'h0000F3A8: begin
				q			<=			16'h0000;
		end
		32'h0000F3AA: begin
				q			<=			16'h0000;
		end
		32'h0000F3AC: begin
				q			<=			16'h9C40;
		end
		32'h0000F3AE: begin
				q			<=			16'h400C;
		end
		32'h0000F3B0: begin
				q			<=			16'h0000;
		end
		32'h0000F3B2: begin
				q			<=			16'h0000;
		end
		32'h0000F3B4: begin
				q			<=			16'h0000;
		end
		32'h0000F3B6: begin
				q			<=			16'h0000;
		end
		32'h0000F3B8: begin
				q			<=			16'h0000;
		end
		32'h0000F3BA: begin
				q			<=			16'h0000;
		end
		32'h0000F3BC: begin
				q			<=			16'h0000;
		end
		32'h0000F3BE: begin
				q			<=			16'h0000;
		end
		32'h0000F3C0: begin
				q			<=			16'hC800;
		end
		32'h0000F3C2: begin
				q			<=			16'h4005;
		end
		32'h0000F3C4: begin
				q			<=			16'h0000;
		end
		32'h0000F3C6: begin
				q			<=			16'h0000;
		end
		32'h0000F3C8: begin
				q			<=			16'h0000;
		end
		32'h0000F3CA: begin
				q			<=			16'h0000;
		end
		32'h0000F3CC: begin
				q			<=			16'h0000;
		end
		32'h0000F3CE: begin
				q			<=			16'h0000;
		end
		32'h0000F3D0: begin
				q			<=			16'h0000;
		end
		32'h0000F3D2: begin
				q			<=			16'h0000;
		end
		32'h0000F3D4: begin
				q			<=			16'hA000;
		end
		32'h0000F3D6: begin
				q			<=			16'h4002;
		end
		32'h0000F3D8: begin
				q			<=			16'hFFFF;
		end
		32'h0000F3DA: begin
				q			<=			16'hFFFE;
		end
		32'h0000F3DC: begin
				q			<=			16'hFFFC;
		end
		32'h0000F3DE: begin
				q			<=			16'hFFF8;
		end
		32'h0000F3E0: begin
				q			<=			16'hFFF0;
		end
		32'h0000F3E2: begin
				q			<=			16'hFFE0;
		end
		32'h0000F3E4: begin
				q			<=			16'hFFC0;
		end
		32'h0000F3E6: begin
				q			<=			16'hFF80;
		end
		32'h0000F3E8: begin
				q			<=			16'hFF00;
		end
		32'h0000F3EA: begin
				q			<=			16'hFE00;
		end
		32'h0000F3EC: begin
				q			<=			16'hFC00;
		end
		32'h0000F3EE: begin
				q			<=			16'hF800;
		end
		32'h0000F3F0: begin
				q			<=			16'hF000;
		end
		32'h0000F3F2: begin
				q			<=			16'hE000;
		end
		32'h0000F3F4: begin
				q			<=			16'hC000;
		end
		32'h0000F3F6: begin
				q			<=			16'h8000;
		end
		32'h0000F3F8: begin
				q			<=			16'h0000;
		end
		32'h0000F3FA: begin
				q			<=			16'h0000;
		end
		32'h0000F3FC: begin
				q			<=			16'h2030;
		end
		32'h0000F3FE: begin
				q			<=			16'hCFFC;
		end
		32'h0000F400: begin
				q			<=			16'hA1C3;
		end
		32'h0000F402: begin
				q			<=			16'h8123;
		end
		32'h0000F404: begin
				q			<=			16'h2DE3;
		end
		32'h0000F406: begin
				q			<=			16'h9FDE;
		end
		32'h0000F408: begin
				q			<=			16'hD2CE;
		end
		32'h0000F40A: begin
				q			<=			16'h04C8;
		end
		32'h0000F40C: begin
				q			<=			16'hA6DD;
		end
		32'h0000F40E: begin
				q			<=			16'h0AD8;
		end
		32'h0000F410: begin
				q			<=			16'h8264;
		end
		32'h0000F412: begin
				q			<=			16'hD2CB;
		end
		32'h0000F414: begin
				q			<=			16'hF2EA;
		end
		32'h0000F416: begin
				q			<=			16'h12D4;
		end
		32'h0000F418: begin
				q			<=			16'h4925;
		end
		32'h0000F41A: begin
				q			<=			16'h2DE4;
		end
		32'h0000F41C: begin
				q			<=			16'h3436;
		end
		32'h0000F41E: begin
				q			<=			16'h534F;
		end
		32'h0000F420: begin
				q			<=			16'hCEAE;
		end
		32'h0000F422: begin
				q			<=			16'h256B;
		end
		32'h0000F424: begin
				q			<=			16'hF53F;
		end
		32'h0000F426: begin
				q			<=			16'hF698;
		end
		32'h0000F428: begin
				q			<=			16'h6BD3;
		end
		32'h0000F42A: begin
				q			<=			16'h0158;
		end
		32'h0000F42C: begin
				q			<=			16'h87A6;
		end
		32'h0000F42E: begin
				q			<=			16'hC0BD;
		end
		32'h0000F430: begin
				q			<=			16'hDA57;
		end
		32'h0000F432: begin
				q			<=			16'h82A5;
		end
		32'h0000F434: begin
				q			<=			16'hA2A6;
		end
		32'h0000F436: begin
				q			<=			16'h32B5;
		end
		32'h0000F438: begin
				q			<=			16'hE731;
		end
		32'h0000F43A: begin
				q			<=			16'h04D4;
		end
		32'h0000F43C: begin
				q			<=			16'hE3F2;
		end
		32'h0000F43E: begin
				q			<=			16'hD332;
		end
		32'h0000F440: begin
				q			<=			16'h7132;
		end
		32'h0000F442: begin
				q			<=			16'hD21C;
		end
		32'h0000F444: begin
				q			<=			16'hDB23;
		end
		32'h0000F446: begin
				q			<=			16'hEE32;
		end
		32'h0000F448: begin
				q			<=			16'h9049;
		end
		32'h0000F44A: begin
				q			<=			16'h395A;
		end
		32'h0000F44C: begin
				q			<=			16'hA23E;
		end
		32'h0000F44E: begin
				q			<=			16'h5308;
		end
		32'h0000F450: begin
				q			<=			16'hFEFB;
		end
		32'h0000F452: begin
				q			<=			16'h1155;
		end
		32'h0000F454: begin
				q			<=			16'hFA91;
		end
		32'h0000F456: begin
				q			<=			16'h1939;
		end
		32'h0000F458: begin
				q			<=			16'h637A;
		end
		32'h0000F45A: begin
				q			<=			16'h4325;
		end
		32'h0000F45C: begin
				q			<=			16'hC031;
		end
		32'h0000F45E: begin
				q			<=			16'h3CAC;
		end
		32'h0000F460: begin
				q			<=			16'hE26D;
		end
		32'h0000F462: begin
				q			<=			16'hDBDE;
		end
		32'h0000F464: begin
				q			<=			16'hD05D;
		end
		32'h0000F466: begin
				q			<=			16'hB3F6;
		end
		32'h0000F468: begin
				q			<=			16'hAC7C;
		end
		32'h0000F46A: begin
				q			<=			16'hE4A0;
		end
		32'h0000F46C: begin
				q			<=			16'h64BC;
		end
		32'h0000F46E: begin
				q			<=			16'h467C;
		end
		32'h0000F470: begin
				q			<=			16'hDDD0;
		end
		32'h0000F472: begin
				q			<=			16'h3E55;
		end
		32'h0000F474: begin
				q			<=			16'h2A20;
		end
		32'h0000F476: begin
				q			<=			16'h6224;
		end
		32'h0000F478: begin
				q			<=			16'h47B3;
		end
		32'h0000F47A: begin
				q			<=			16'h98D7;
		end
		32'h0000F47C: begin
				q			<=			16'h3F23;
		end
		32'h0000F47E: begin
				q			<=			16'hE9A5;
		end
		32'h0000F480: begin
				q			<=			16'hA539;
		end
		32'h0000F482: begin
				q			<=			16'hEA27;
		end
		32'h0000F484: begin
				q			<=			16'hA87F;
		end
		32'h0000F486: begin
				q			<=			16'h3F2A;
		end
		32'h0000F488: begin
				q			<=			16'h0B5B;
		end
		32'h0000F48A: begin
				q			<=			16'h4AF2;
		end
		32'h0000F48C: begin
				q			<=			16'hA581;
		end
		32'h0000F48E: begin
				q			<=			16'h18ED;
		end
		32'h0000F490: begin
				q			<=			16'h67DE;
		end
		32'h0000F492: begin
				q			<=			16'h94BA;
		end
		32'h0000F494: begin
				q			<=			16'h4539;
		end
		32'h0000F496: begin
				q			<=			16'h1EAD;
		end
		32'h0000F498: begin
				q			<=			16'hCFB1;
		end
		32'h0000F49A: begin
				q			<=			16'h3F94;
		end
		32'h0000F49C: begin
				q			<=			16'hBF71;
		end
		32'h0000F49E: begin
				q			<=			16'hA9B3;
		end
		32'h0000F4A0: begin
				q			<=			16'h7989;
		end
		32'h0000F4A2: begin
				q			<=			16'hBE68;
		end
		32'h0000F4A4: begin
				q			<=			16'h4C2E;
		end
		32'h0000F4A6: begin
				q			<=			16'hE15B;
		end
		32'h0000F4A8: begin
				q			<=			16'hC44D;
		end
		32'h0000F4AA: begin
				q			<=			16'h94BE;
		end
		32'h0000F4AC: begin
				q			<=			16'hE695;
		end
		32'h0000F4AE: begin
				q			<=			16'h3FC9;
		end
		32'h0000F4B0: begin
				q			<=			16'h3D4D;
		end
		32'h0000F4B2: begin
				q			<=			16'h7C3D;
		end
		32'h0000F4B4: begin
				q			<=			16'h36BA;
		end
		32'h0000F4B6: begin
				q			<=			16'h0D2B;
		end
		32'h0000F4B8: begin
				q			<=			16'hFDC2;
		end
		32'h0000F4BA: begin
				q			<=			16'hCEFC;
		end
		32'h0000F4BC: begin
				q			<=			16'h8461;
		end
		32'h0000F4BE: begin
				q			<=			16'h7711;
		end
		32'h0000F4C0: begin
				q			<=			16'hABCC;
		end
		32'h0000F4C2: begin
				q			<=			16'h3FE4;
		end
		32'h0000F4C4: begin
				q			<=			16'hC155;
		end
		32'h0000F4C6: begin
				q			<=			16'hA4A8;
		end
		32'h0000F4C8: begin
				q			<=			16'h404E;
		end
		32'h0000F4CA: begin
				q			<=			16'h6113;
		end
		32'h0000F4CC: begin
				q			<=			16'hD3C3;
		end
		32'h0000F4CE: begin
				q			<=			16'h652B;
		end
		32'h0000F4D0: begin
				q			<=			16'hE219;
		end
		32'h0000F4D2: begin
				q			<=			16'h1758;
		end
		32'h0000F4D4: begin
				q			<=			16'hD1B7;
		end
		32'h0000F4D6: begin
				q			<=			16'h3FF1;
		end
		32'h0000F4D8: begin
				q			<=			16'hD70A;
		end
		32'h0000F4DA: begin
				q			<=			16'h70A3;
		end
		32'h0000F4DC: begin
				q			<=			16'h0A3D;
		end
		32'h0000F4DE: begin
				q			<=			16'hA3D7;
		end
		32'h0000F4E0: begin
				q			<=			16'h3D70;
		end
		32'h0000F4E2: begin
				q			<=			16'hD70A;
		end
		32'h0000F4E4: begin
				q			<=			16'h70A3;
		end
		32'h0000F4E6: begin
				q			<=			16'h0A3D;
		end
		32'h0000F4E8: begin
				q			<=			16'hA3D7;
		end
		32'h0000F4EA: begin
				q			<=			16'h3FF8;
		end
		32'h0000F4EC: begin
				q			<=			16'hCCCD;
		end
		32'h0000F4EE: begin
				q			<=			16'hCCCC;
		end
		32'h0000F4F0: begin
				q			<=			16'hCCCC;
		end
		32'h0000F4F2: begin
				q			<=			16'hCCCC;
		end
		32'h0000F4F4: begin
				q			<=			16'hCCCC;
		end
		32'h0000F4F6: begin
				q			<=			16'hCCCC;
		end
		32'h0000F4F8: begin
				q			<=			16'hCCCC;
		end
		32'h0000F4FA: begin
				q			<=			16'hCCCC;
		end
		32'h0000F4FC: begin
				q			<=			16'hCCCC;
		end
		32'h0000F4FE: begin
				q			<=			16'h3FFB;
		end
		32'h0000F500: begin
				q			<=			16'h0005;
		end
		32'h0000F502: begin
				q			<=			16'h0000;
		end
		32'h0000F504: begin
				q			<=			16'h0019;
		end
		32'h0000F506: begin
				q			<=			16'h0000;
		end
		32'h0000F508: begin
				q			<=			16'h007D;
		end
		32'h0000F50A: begin
				q			<=			16'h0000;
		end
		32'h0000F50C: begin
				q			<=			16'h0000;
		end
		32'h0000F50E: begin
				q			<=			16'h0000;
		end
		32'h0000F510: begin
				q			<=			16'h0000;
		end
		32'h0000F512: begin
				q			<=			16'h0000;
		end
		32'h0000F514: begin
				q			<=			16'h0000;
		end
		32'h0000F516: begin
				q			<=			16'h3FF0;
		end
		32'h0000F518: begin
				q			<=			16'h0000;
		end
		32'h0000F51A: begin
				q			<=			16'h0000;
		end
		32'h0000F51C: begin
				q			<=			16'h0000;
		end
		32'h0000F51E: begin
				q			<=			16'h4024;
		end
		32'h0000F520: begin
				q			<=			16'h0000;
		end
		32'h0000F522: begin
				q			<=			16'h0000;
		end
		32'h0000F524: begin
				q			<=			16'h0000;
		end
		32'h0000F526: begin
				q			<=			16'h4059;
		end
		32'h0000F528: begin
				q			<=			16'h0000;
		end
		32'h0000F52A: begin
				q			<=			16'h0000;
		end
		32'h0000F52C: begin
				q			<=			16'h4000;
		end
		32'h0000F52E: begin
				q			<=			16'h408F;
		end
		32'h0000F530: begin
				q			<=			16'h0000;
		end
		32'h0000F532: begin
				q			<=			16'h0000;
		end
		32'h0000F534: begin
				q			<=			16'h8800;
		end
		32'h0000F536: begin
				q			<=			16'h40C3;
		end
		32'h0000F538: begin
				q			<=			16'h0000;
		end
		32'h0000F53A: begin
				q			<=			16'h0000;
		end
		32'h0000F53C: begin
				q			<=			16'h6A00;
		end
		32'h0000F53E: begin
				q			<=			16'h40F8;
		end
		32'h0000F540: begin
				q			<=			16'h0000;
		end
		32'h0000F542: begin
				q			<=			16'h0000;
		end
		32'h0000F544: begin
				q			<=			16'h8480;
		end
		32'h0000F546: begin
				q			<=			16'h412E;
		end
		32'h0000F548: begin
				q			<=			16'h0000;
		end
		32'h0000F54A: begin
				q			<=			16'h0000;
		end
		32'h0000F54C: begin
				q			<=			16'h12D0;
		end
		32'h0000F54E: begin
				q			<=			16'h4163;
		end
		32'h0000F550: begin
				q			<=			16'h0000;
		end
		32'h0000F552: begin
				q			<=			16'h0000;
		end
		32'h0000F554: begin
				q			<=			16'hD784;
		end
		32'h0000F556: begin
				q			<=			16'h4197;
		end
		32'h0000F558: begin
				q			<=			16'h0000;
		end
		32'h0000F55A: begin
				q			<=			16'h0000;
		end
		32'h0000F55C: begin
				q			<=			16'hCD65;
		end
		32'h0000F55E: begin
				q			<=			16'h41CD;
		end
		32'h0000F560: begin
				q			<=			16'h0000;
		end
		32'h0000F562: begin
				q			<=			16'h2000;
		end
		32'h0000F564: begin
				q			<=			16'hA05F;
		end
		32'h0000F566: begin
				q			<=			16'h4202;
		end
		32'h0000F568: begin
				q			<=			16'h0000;
		end
		32'h0000F56A: begin
				q			<=			16'hE800;
		end
		32'h0000F56C: begin
				q			<=			16'h4876;
		end
		32'h0000F56E: begin
				q			<=			16'h4237;
		end
		32'h0000F570: begin
				q			<=			16'h0000;
		end
		32'h0000F572: begin
				q			<=			16'hA200;
		end
		32'h0000F574: begin
				q			<=			16'h1A94;
		end
		32'h0000F576: begin
				q			<=			16'h426D;
		end
		32'h0000F578: begin
				q			<=			16'h0000;
		end
		32'h0000F57A: begin
				q			<=			16'hE540;
		end
		32'h0000F57C: begin
				q			<=			16'h309C;
		end
		32'h0000F57E: begin
				q			<=			16'h42A2;
		end
		32'h0000F580: begin
				q			<=			16'h0000;
		end
		32'h0000F582: begin
				q			<=			16'h1E90;
		end
		32'h0000F584: begin
				q			<=			16'hBCC4;
		end
		32'h0000F586: begin
				q			<=			16'h42D6;
		end
		32'h0000F588: begin
				q			<=			16'h0000;
		end
		32'h0000F58A: begin
				q			<=			16'h2634;
		end
		32'h0000F58C: begin
				q			<=			16'h6BF5;
		end
		32'h0000F58E: begin
				q			<=			16'h430C;
		end
		32'h0000F590: begin
				q			<=			16'h8000;
		end
		32'h0000F592: begin
				q			<=			16'h37E0;
		end
		32'h0000F594: begin
				q			<=			16'hC379;
		end
		32'h0000F596: begin
				q			<=			16'h4341;
		end
		32'h0000F598: begin
				q			<=			16'hA000;
		end
		32'h0000F59A: begin
				q			<=			16'h85D8;
		end
		32'h0000F59C: begin
				q			<=			16'h3457;
		end
		32'h0000F59E: begin
				q			<=			16'h4376;
		end
		32'h0000F5A0: begin
				q			<=			16'hC800;
		end
		32'h0000F5A2: begin
				q			<=			16'h674E;
		end
		32'h0000F5A4: begin
				q			<=			16'hC16D;
		end
		32'h0000F5A6: begin
				q			<=			16'h43AB;
		end
		32'h0000F5A8: begin
				q			<=			16'h3D00;
		end
		32'h0000F5AA: begin
				q			<=			16'h6091;
		end
		32'h0000F5AC: begin
				q			<=			16'h58E4;
		end
		32'h0000F5AE: begin
				q			<=			16'h43E1;
		end
		32'h0000F5B0: begin
				q			<=			16'h8C40;
		end
		32'h0000F5B2: begin
				q			<=			16'h78B5;
		end
		32'h0000F5B4: begin
				q			<=			16'hAF1D;
		end
		32'h0000F5B6: begin
				q			<=			16'h4415;
		end
		32'h0000F5B8: begin
				q			<=			16'hEF50;
		end
		32'h0000F5BA: begin
				q			<=			16'hD6E2;
		end
		32'h0000F5BC: begin
				q			<=			16'h1AE4;
		end
		32'h0000F5BE: begin
				q			<=			16'h444B;
		end
		32'h0000F5C0: begin
				q			<=			16'hD592;
		end
		32'h0000F5C2: begin
				q			<=			16'h064D;
		end
		32'h0000F5C4: begin
				q			<=			16'hF0CF;
		end
		32'h0000F5C6: begin
				q			<=			16'h4480;
		end
		32'h0000F5C8: begin
				q			<=			16'h4AF6;
		end
		32'h0000F5CA: begin
				q			<=			16'hC7E1;
		end
		32'h0000F5CC: begin
				q			<=			16'h2D02;
		end
		32'h0000F5CE: begin
				q			<=			16'h44B5;
		end
		32'h0000F5D0: begin
				q			<=			16'h9DB4;
		end
		32'h0000F5D2: begin
				q			<=			16'h79D9;
		end
		32'h0000F5D4: begin
				q			<=			16'h7843;
		end
		32'h0000F5D6: begin
				q			<=			16'h44EA;
		end
		32'h0000F5D8: begin
				q			<=			16'h89BC;
		end
		32'h0000F5DA: begin
				q			<=			16'h97D8;
		end
		32'h0000F5DC: begin
				q			<=			16'hD2B2;
		end
		32'h0000F5DE: begin
				q			<=			16'h3C9C;
		end
		32'h0000F5E0: begin
				q			<=			16'hA733;
		end
		32'h0000F5E2: begin
				q			<=			16'hD5A8;
		end
		32'h0000F5E4: begin
				q			<=			16'hF623;
		end
		32'h0000F5E6: begin
				q			<=			16'h3949;
		end
		32'h0000F5E8: begin
				q			<=			16'hA73D;
		end
		32'h0000F5EA: begin
				q			<=			16'h44F4;
		end
		32'h0000F5EC: begin
				q			<=			16'h0FFD;
		end
		32'h0000F5EE: begin
				q			<=			16'h32A5;
		end
		32'h0000F5F0: begin
				q			<=			16'h979D;
		end
		32'h0000F5F2: begin
				q			<=			16'hCF8C;
		end
		32'h0000F5F4: begin
				q			<=			16'hBA08;
		end
		32'h0000F5F6: begin
				q			<=			16'h255B;
		end
		32'h0000F5F8: begin
				q			<=			16'h6F43;
		end
		32'h0000F5FA: begin
				q			<=			16'h64AC;
		end
		32'h0000F5FC: begin
				q			<=			16'h0628;
		end
		32'h0000F5FE: begin
				q			<=			16'h0AC8;
		end
		32'h0000F600: begin
				q			<=			16'h8000;
		end
		32'h0000F602: begin
				q			<=			16'h37E0;
		end
		32'h0000F604: begin
				q			<=			16'hC379;
		end
		32'h0000F606: begin
				q			<=			16'h4341;
		end
		32'h0000F608: begin
				q			<=			16'h6E17;
		end
		32'h0000F60A: begin
				q			<=			16'hB505;
		end
		32'h0000F60C: begin
				q			<=			16'hB8B5;
		end
		32'h0000F60E: begin
				q			<=			16'h4693;
		end
		32'h0000F610: begin
				q			<=			16'hF9F5;
		end
		32'h0000F612: begin
				q			<=			16'hE93F;
		end
		32'h0000F614: begin
				q			<=			16'h4F03;
		end
		32'h0000F616: begin
				q			<=			16'h4D38;
		end
		32'h0000F618: begin
				q			<=			16'h1D32;
		end
		32'h0000F61A: begin
				q			<=			16'hF930;
		end
		32'h0000F61C: begin
				q			<=			16'h7748;
		end
		32'h0000F61E: begin
				q			<=			16'h5A82;
		end
		32'h0000F620: begin
				q			<=			16'hBF3C;
		end
		32'h0000F622: begin
				q			<=			16'h7F73;
		end
		32'h0000F624: begin
				q			<=			16'h4FDD;
		end
		32'h0000F626: begin
				q			<=			16'h7515;
		end
		32'h0000F628: begin
				q			<=			16'h9920;
		end
		32'h0000F62A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F62C: begin
				q			<=			16'hA178;
		end
		32'h0000F62E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F630: begin
				q			<=			16'hA178;
		end
		32'h0000F632: begin
				q			<=			16'hFFFF;
		end
		32'h0000F634: begin
				q			<=			16'h9934;
		end
		32'h0000F636: begin
				q			<=			16'hFFFF;
		end
		32'h0000F638: begin
				q			<=			16'hA178;
		end
		32'h0000F63A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F63C: begin
				q			<=			16'hA178;
		end
		32'h0000F63E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F640: begin
				q			<=			16'hA178;
		end
		32'h0000F642: begin
				q			<=			16'hFFFF;
		end
		32'h0000F644: begin
				q			<=			16'h98C8;
		end
		32'h0000F646: begin
				q			<=			16'hFFFF;
		end
		32'h0000F648: begin
				q			<=			16'hA178;
		end
		32'h0000F64A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F64C: begin
				q			<=			16'hA178;
		end
		32'h0000F64E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F650: begin
				q			<=			16'h993C;
		end
		32'h0000F652: begin
				q			<=			16'hFFFF;
		end
		32'h0000F654: begin
				q			<=			16'h9954;
		end
		32'h0000F656: begin
				q			<=			16'hFFFF;
		end
		32'h0000F658: begin
				q			<=			16'hA178;
		end
		32'h0000F65A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F65C: begin
				q			<=			16'h994C;
		end
		32'h0000F65E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F660: begin
				q			<=			16'h995C;
		end
		32'h0000F662: begin
				q			<=			16'hFFFF;
		end
		32'h0000F664: begin
				q			<=			16'hA178;
		end
		32'h0000F666: begin
				q			<=			16'hFFFF;
		end
		32'h0000F668: begin
				q			<=			16'h99B0;
		end
		32'h0000F66A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F66C: begin
				q			<=			16'h99B8;
		end
		32'h0000F66E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F670: begin
				q			<=			16'h99B8;
		end
		32'h0000F672: begin
				q			<=			16'hFFFF;
		end
		32'h0000F674: begin
				q			<=			16'h99B8;
		end
		32'h0000F676: begin
				q			<=			16'hFFFF;
		end
		32'h0000F678: begin
				q			<=			16'h99B8;
		end
		32'h0000F67A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F67C: begin
				q			<=			16'h99B8;
		end
		32'h0000F67E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F680: begin
				q			<=			16'h99B8;
		end
		32'h0000F682: begin
				q			<=			16'hFFFF;
		end
		32'h0000F684: begin
				q			<=			16'h99B8;
		end
		32'h0000F686: begin
				q			<=			16'hFFFF;
		end
		32'h0000F688: begin
				q			<=			16'h99B8;
		end
		32'h0000F68A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F68C: begin
				q			<=			16'h99B8;
		end
		32'h0000F68E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F690: begin
				q			<=			16'hA178;
		end
		32'h0000F692: begin
				q			<=			16'hFFFF;
		end
		32'h0000F694: begin
				q			<=			16'hA178;
		end
		32'h0000F696: begin
				q			<=			16'hFFFF;
		end
		32'h0000F698: begin
				q			<=			16'hA178;
		end
		32'h0000F69A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F69C: begin
				q			<=			16'hA178;
		end
		32'h0000F69E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6A0: begin
				q			<=			16'hA178;
		end
		32'h0000F6A2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6A4: begin
				q			<=			16'hA178;
		end
		32'h0000F6A6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6A8: begin
				q			<=			16'hA178;
		end
		32'h0000F6AA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6AC: begin
				q			<=			16'hA178;
		end
		32'h0000F6AE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6B0: begin
				q			<=			16'hA178;
		end
		32'h0000F6B2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6B4: begin
				q			<=			16'h9A24;
		end
		32'h0000F6B6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6B8: begin
				q			<=			16'h9A44;
		end
		32'h0000F6BA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6BC: begin
				q			<=			16'hA178;
		end
		32'h0000F6BE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6C0: begin
				q			<=			16'hA178;
		end
		32'h0000F6C2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6C4: begin
				q			<=			16'hA178;
		end
		32'h0000F6C6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6C8: begin
				q			<=			16'hA178;
		end
		32'h0000F6CA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6CC: begin
				q			<=			16'hA178;
		end
		32'h0000F6CE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6D0: begin
				q			<=			16'hA178;
		end
		32'h0000F6D2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6D4: begin
				q			<=			16'hA178;
		end
		32'h0000F6D6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6D8: begin
				q			<=			16'hA178;
		end
		32'h0000F6DA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6DC: begin
				q			<=			16'hA178;
		end
		32'h0000F6DE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6E0: begin
				q			<=			16'hA178;
		end
		32'h0000F6E2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6E4: begin
				q			<=			16'h9B38;
		end
		32'h0000F6E6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6E8: begin
				q			<=			16'hA178;
		end
		32'h0000F6EA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6EC: begin
				q			<=			16'hA178;
		end
		32'h0000F6EE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6F0: begin
				q			<=			16'hA178;
		end
		32'h0000F6F2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6F4: begin
				q			<=			16'h9BF4;
		end
		32'h0000F6F6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6F8: begin
				q			<=			16'hA178;
		end
		32'h0000F6FA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F6FC: begin
				q			<=			16'h9F14;
		end
		32'h0000F6FE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F700: begin
				q			<=			16'hA178;
		end
		32'h0000F702: begin
				q			<=			16'hFFFF;
		end
		32'h0000F704: begin
				q			<=			16'hA178;
		end
		32'h0000F706: begin
				q			<=			16'hFFFF;
		end
		32'h0000F708: begin
				q			<=			16'h9878;
		end
		32'h0000F70A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F70C: begin
				q			<=			16'hA178;
		end
		32'h0000F70E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F710: begin
				q			<=			16'hA178;
		end
		32'h0000F712: begin
				q			<=			16'hFFFF;
		end
		32'h0000F714: begin
				q			<=			16'hA178;
		end
		32'h0000F716: begin
				q			<=			16'hFFFF;
		end
		32'h0000F718: begin
				q			<=			16'hA178;
		end
		32'h0000F71A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F71C: begin
				q			<=			16'hA178;
		end
		32'h0000F71E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F720: begin
				q			<=			16'hA178;
		end
		32'h0000F722: begin
				q			<=			16'hFFFF;
		end
		32'h0000F724: begin
				q			<=			16'hA178;
		end
		32'h0000F726: begin
				q			<=			16'hFFFF;
		end
		32'h0000F728: begin
				q			<=			16'hA178;
		end
		32'h0000F72A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F72C: begin
				q			<=			16'hA178;
		end
		32'h0000F72E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F730: begin
				q			<=			16'hA178;
		end
		32'h0000F732: begin
				q			<=			16'hFFFF;
		end
		32'h0000F734: begin
				q			<=			16'h9A24;
		end
		32'h0000F736: begin
				q			<=			16'hFFFF;
		end
		32'h0000F738: begin
				q			<=			16'h9A48;
		end
		32'h0000F73A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F73C: begin
				q			<=			16'hA178;
		end
		32'h0000F73E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F740: begin
				q			<=			16'hA178;
		end
		32'h0000F742: begin
				q			<=			16'hFFFF;
		end
		32'h0000F744: begin
				q			<=			16'hA178;
		end
		32'h0000F746: begin
				q			<=			16'hFFFF;
		end
		32'h0000F748: begin
				q			<=			16'h99E4;
		end
		32'h0000F74A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F74C: begin
				q			<=			16'h9A48;
		end
		32'h0000F74E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F750: begin
				q			<=			16'h9A14;
		end
		32'h0000F752: begin
				q			<=			16'hFFFF;
		end
		32'h0000F754: begin
				q			<=			16'hA178;
		end
		32'h0000F756: begin
				q			<=			16'hFFFF;
		end
		32'h0000F758: begin
				q			<=			16'h9A04;
		end
		32'h0000F75A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F75C: begin
				q			<=			16'hA178;
		end
		32'h0000F75E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F760: begin
				q			<=			16'h9AE8;
		end
		32'h0000F762: begin
				q			<=			16'hFFFF;
		end
		32'h0000F764: begin
				q			<=			16'h9B3C;
		end
		32'h0000F766: begin
				q			<=			16'hFFFF;
		end
		32'h0000F768: begin
				q			<=			16'h9BC4;
		end
		32'h0000F76A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F76C: begin
				q			<=			16'h9A14;
		end
		32'h0000F76E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F770: begin
				q			<=			16'hA178;
		end
		32'h0000F772: begin
				q			<=			16'hFFFF;
		end
		32'h0000F774: begin
				q			<=			16'h9BF4;
		end
		32'h0000F776: begin
				q			<=			16'hFFFF;
		end
		32'h0000F778: begin
				q			<=			16'h9844;
		end
		32'h0000F77A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F77C: begin
				q			<=			16'h9F18;
		end
		32'h0000F77E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F780: begin
				q			<=			16'hA178;
		end
		32'h0000F782: begin
				q			<=			16'hFFFF;
		end
		32'h0000F784: begin
				q			<=			16'hA178;
		end
		32'h0000F786: begin
				q			<=			16'hFFFF;
		end
		32'h0000F788: begin
				q			<=			16'h9F74;
		end
		32'h0000F78A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F78C: begin
				q			<=			16'hA178;
		end
		32'h0000F78E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F790: begin
				q			<=			16'h9844;
		end
		32'h0000F792: begin
				q			<=			16'hFFFF;
		end
		32'h0000F794: begin
				q			<=			16'h2020;
		end
		32'h0000F796: begin
				q			<=			16'h2020;
		end
		32'h0000F798: begin
				q			<=			16'h2020;
		end
		32'h0000F79A: begin
				q			<=			16'h2020;
		end
		32'h0000F79C: begin
				q			<=			16'h2020;
		end
		32'h0000F79E: begin
				q			<=			16'h2020;
		end
		32'h0000F7A0: begin
				q			<=			16'h2020;
		end
		32'h0000F7A2: begin
				q			<=			16'h2020;
		end
		32'h0000F7A4: begin
				q			<=			16'h3030;
		end
		32'h0000F7A6: begin
				q			<=			16'h3030;
		end
		32'h0000F7A8: begin
				q			<=			16'h3030;
		end
		32'h0000F7AA: begin
				q			<=			16'h3030;
		end
		32'h0000F7AC: begin
				q			<=			16'h3030;
		end
		32'h0000F7AE: begin
				q			<=			16'h3030;
		end
		32'h0000F7B0: begin
				q			<=			16'h3030;
		end
		32'h0000F7B2: begin
				q			<=			16'h3030;
		end
		32'h0000F7B4: begin
				q			<=			16'h2000;
		end
		32'h0000F7B6: begin
				q			<=			16'h2020;
		end
		32'h0000F7B8: begin
				q			<=			16'h2020;
		end
		32'h0000F7BA: begin
				q			<=			16'h2020;
		end
		32'h0000F7BC: begin
				q			<=			16'h2020;
		end
		32'h0000F7BE: begin
				q			<=			16'h2828;
		end
		32'h0000F7C0: begin
				q			<=			16'h2828;
		end
		32'h0000F7C2: begin
				q			<=			16'h2028;
		end
		32'h0000F7C4: begin
				q			<=			16'h2020;
		end
		32'h0000F7C6: begin
				q			<=			16'h2020;
		end
		32'h0000F7C8: begin
				q			<=			16'h2020;
		end
		32'h0000F7CA: begin
				q			<=			16'h2020;
		end
		32'h0000F7CC: begin
				q			<=			16'h2020;
		end
		32'h0000F7CE: begin
				q			<=			16'h2020;
		end
		32'h0000F7D0: begin
				q			<=			16'h2020;
		end
		32'h0000F7D2: begin
				q			<=			16'h2020;
		end
		32'h0000F7D4: begin
				q			<=			16'h8820;
		end
		32'h0000F7D6: begin
				q			<=			16'h1010;
		end
		32'h0000F7D8: begin
				q			<=			16'h1010;
		end
		32'h0000F7DA: begin
				q			<=			16'h1010;
		end
		32'h0000F7DC: begin
				q			<=			16'h1010;
		end
		32'h0000F7DE: begin
				q			<=			16'h1010;
		end
		32'h0000F7E0: begin
				q			<=			16'h1010;
		end
		32'h0000F7E2: begin
				q			<=			16'h1010;
		end
		32'h0000F7E4: begin
				q			<=			16'h0410;
		end
		32'h0000F7E6: begin
				q			<=			16'h0404;
		end
		32'h0000F7E8: begin
				q			<=			16'h0404;
		end
		32'h0000F7EA: begin
				q			<=			16'h0404;
		end
		32'h0000F7EC: begin
				q			<=			16'h0404;
		end
		32'h0000F7EE: begin
				q			<=			16'h1004;
		end
		32'h0000F7F0: begin
				q			<=			16'h1010;
		end
		32'h0000F7F2: begin
				q			<=			16'h1010;
		end
		32'h0000F7F4: begin
				q			<=			16'h1010;
		end
		32'h0000F7F6: begin
				q			<=			16'h4141;
		end
		32'h0000F7F8: begin
				q			<=			16'h4141;
		end
		32'h0000F7FA: begin
				q			<=			16'h4141;
		end
		32'h0000F7FC: begin
				q			<=			16'h0101;
		end
		32'h0000F7FE: begin
				q			<=			16'h0101;
		end
		32'h0000F800: begin
				q			<=			16'h0101;
		end
		32'h0000F802: begin
				q			<=			16'h0101;
		end
		32'h0000F804: begin
				q			<=			16'h0101;
		end
		32'h0000F806: begin
				q			<=			16'h0101;
		end
		32'h0000F808: begin
				q			<=			16'h0101;
		end
		32'h0000F80A: begin
				q			<=			16'h0101;
		end
		32'h0000F80C: begin
				q			<=			16'h0101;
		end
		32'h0000F80E: begin
				q			<=			16'h0101;
		end
		32'h0000F810: begin
				q			<=			16'h1010;
		end
		32'h0000F812: begin
				q			<=			16'h1010;
		end
		32'h0000F814: begin
				q			<=			16'h1010;
		end
		32'h0000F816: begin
				q			<=			16'h4242;
		end
		32'h0000F818: begin
				q			<=			16'h4242;
		end
		32'h0000F81A: begin
				q			<=			16'h4242;
		end
		32'h0000F81C: begin
				q			<=			16'h0202;
		end
		32'h0000F81E: begin
				q			<=			16'h0202;
		end
		32'h0000F820: begin
				q			<=			16'h0202;
		end
		32'h0000F822: begin
				q			<=			16'h0202;
		end
		32'h0000F824: begin
				q			<=			16'h0202;
		end
		32'h0000F826: begin
				q			<=			16'h0202;
		end
		32'h0000F828: begin
				q			<=			16'h0202;
		end
		32'h0000F82A: begin
				q			<=			16'h0202;
		end
		32'h0000F82C: begin
				q			<=			16'h0202;
		end
		32'h0000F82E: begin
				q			<=			16'h0202;
		end
		32'h0000F830: begin
				q			<=			16'h1010;
		end
		32'h0000F832: begin
				q			<=			16'h1010;
		end
		32'h0000F834: begin
				q			<=			16'h0020;
		end
		32'h0000F836: begin
				q			<=			16'h0000;
		end
		32'h0000F838: begin
				q			<=			16'h0000;
		end
		32'h0000F83A: begin
				q			<=			16'h0000;
		end
		32'h0000F83C: begin
				q			<=			16'h0000;
		end
		32'h0000F83E: begin
				q			<=			16'h0000;
		end
		32'h0000F840: begin
				q			<=			16'h0000;
		end
		32'h0000F842: begin
				q			<=			16'h0000;
		end
		32'h0000F844: begin
				q			<=			16'h0000;
		end
		32'h0000F846: begin
				q			<=			16'h0000;
		end
		32'h0000F848: begin
				q			<=			16'h0000;
		end
		32'h0000F84A: begin
				q			<=			16'h0000;
		end
		32'h0000F84C: begin
				q			<=			16'h0000;
		end
		32'h0000F84E: begin
				q			<=			16'h0000;
		end
		32'h0000F850: begin
				q			<=			16'h0000;
		end
		32'h0000F852: begin
				q			<=			16'h0000;
		end
		32'h0000F854: begin
				q			<=			16'h0000;
		end
		32'h0000F856: begin
				q			<=			16'h0000;
		end
		32'h0000F858: begin
				q			<=			16'h0000;
		end
		32'h0000F85A: begin
				q			<=			16'h0000;
		end
		32'h0000F85C: begin
				q			<=			16'h0000;
		end
		32'h0000F85E: begin
				q			<=			16'h0000;
		end
		32'h0000F860: begin
				q			<=			16'h0000;
		end
		32'h0000F862: begin
				q			<=			16'h0000;
		end
		32'h0000F864: begin
				q			<=			16'h0000;
		end
		32'h0000F866: begin
				q			<=			16'h0000;
		end
		32'h0000F868: begin
				q			<=			16'h0000;
		end
		32'h0000F86A: begin
				q			<=			16'h0000;
		end
		32'h0000F86C: begin
				q			<=			16'h0000;
		end
		32'h0000F86E: begin
				q			<=			16'h0000;
		end
		32'h0000F870: begin
				q			<=			16'h0000;
		end
		32'h0000F872: begin
				q			<=			16'h0000;
		end
		32'h0000F874: begin
				q			<=			16'h0000;
		end
		32'h0000F876: begin
				q			<=			16'h0000;
		end
		32'h0000F878: begin
				q			<=			16'h0000;
		end
		32'h0000F87A: begin
				q			<=			16'h0000;
		end
		32'h0000F87C: begin
				q			<=			16'h0000;
		end
		32'h0000F87E: begin
				q			<=			16'h0000;
		end
		32'h0000F880: begin
				q			<=			16'h0000;
		end
		32'h0000F882: begin
				q			<=			16'h0000;
		end
		32'h0000F884: begin
				q			<=			16'h0000;
		end
		32'h0000F886: begin
				q			<=			16'h0000;
		end
		32'h0000F888: begin
				q			<=			16'h0000;
		end
		32'h0000F88A: begin
				q			<=			16'h0000;
		end
		32'h0000F88C: begin
				q			<=			16'h0000;
		end
		32'h0000F88E: begin
				q			<=			16'h0000;
		end
		32'h0000F890: begin
				q			<=			16'h0000;
		end
		32'h0000F892: begin
				q			<=			16'h0000;
		end
		32'h0000F894: begin
				q			<=			16'h0000;
		end
		32'h0000F896: begin
				q			<=			16'h0000;
		end
		32'h0000F898: begin
				q			<=			16'h0000;
		end
		32'h0000F89A: begin
				q			<=			16'h0000;
		end
		32'h0000F89C: begin
				q			<=			16'h0000;
		end
		32'h0000F89E: begin
				q			<=			16'h0000;
		end
		32'h0000F8A0: begin
				q			<=			16'h0000;
		end
		32'h0000F8A2: begin
				q			<=			16'h0000;
		end
		32'h0000F8A4: begin
				q			<=			16'h0000;
		end
		32'h0000F8A6: begin
				q			<=			16'h0000;
		end
		32'h0000F8A8: begin
				q			<=			16'h0000;
		end
		32'h0000F8AA: begin
				q			<=			16'h0000;
		end
		32'h0000F8AC: begin
				q			<=			16'h0000;
		end
		32'h0000F8AE: begin
				q			<=			16'h0000;
		end
		32'h0000F8B0: begin
				q			<=			16'h0000;
		end
		32'h0000F8B2: begin
				q			<=			16'h0000;
		end
		32'h0000F8B4: begin
				q			<=			16'h0000;
		end
		32'h0000F8B6: begin
				q			<=			16'h0000;
		end
		32'h0000F8B8: begin
				q			<=			16'hC100;
		end
		32'h0000F8BA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8BC: begin
				q			<=			16'hC014;
		end
		32'h0000F8BE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8C0: begin
				q			<=			16'hC020;
		end
		32'h0000F8C2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8C4: begin
				q			<=			16'hC014;
		end
		32'h0000F8C6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8C8: begin
				q			<=			16'hC0EC;
		end
		32'h0000F8CA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8CC: begin
				q			<=			16'hC014;
		end
		32'h0000F8CE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8D0: begin
				q			<=			16'hC020;
		end
		32'h0000F8D2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8D4: begin
				q			<=			16'hC100;
		end
		32'h0000F8D6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8D8: begin
				q			<=			16'hC100;
		end
		32'h0000F8DA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8DC: begin
				q			<=			16'hC0EC;
		end
		32'h0000F8DE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8E0: begin
				q			<=			16'hC020;
		end
		32'h0000F8E2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8E4: begin
				q			<=			16'hBFEC;
		end
		32'h0000F8E6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8E8: begin
				q			<=			16'hBFEC;
		end
		32'h0000F8EA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8EC: begin
				q			<=			16'hBFEC;
		end
		32'h0000F8EE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8F0: begin
				q			<=			16'hC028;
		end
		32'h0000F8F2: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8F4: begin
				q			<=			16'hC5AC;
		end
		32'h0000F8F6: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8F8: begin
				q			<=			16'hC5AC;
		end
		32'h0000F8FA: begin
				q			<=			16'hFFFF;
		end
		32'h0000F8FC: begin
				q			<=			16'hC5D0;
		end
		32'h0000F8FE: begin
				q			<=			16'hFFFF;
		end
		32'h0000F900: begin
				q			<=			16'hC5A0;
		end
		32'h0000F902: begin
				q			<=			16'hFFFF;
		end
		32'h0000F904: begin
				q			<=			16'hC5A0;
		end
		32'h0000F906: begin
				q			<=			16'hFFFF;
		end
		32'h0000F908: begin
				q			<=			16'hC690;
		end
		32'h0000F90A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F90C: begin
				q			<=			16'hC5D0;
		end
		32'h0000F90E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F910: begin
				q			<=			16'hC5A0;
		end
		32'h0000F912: begin
				q			<=			16'hFFFF;
		end
		32'h0000F914: begin
				q			<=			16'hC690;
		end
		32'h0000F916: begin
				q			<=			16'hFFFF;
		end
		32'h0000F918: begin
				q			<=			16'hC5A0;
		end
		32'h0000F91A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F91C: begin
				q			<=			16'hC5D0;
		end
		32'h0000F91E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F920: begin
				q			<=			16'hC59C;
		end
		32'h0000F922: begin
				q			<=			16'hFFFF;
		end
		32'h0000F924: begin
				q			<=			16'hC59C;
		end
		32'h0000F926: begin
				q			<=			16'hFFFF;
		end
		32'h0000F928: begin
				q			<=			16'hC59C;
		end
		32'h0000F92A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F92C: begin
				q			<=			16'hC690;
		end
		32'h0000F92E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F930: begin
				q			<=			16'hD7D4;
		end
		32'h0000F932: begin
				q			<=			16'hFFFF;
		end
		32'h0000F934: begin
				q			<=			16'hD7D4;
		end
		32'h0000F936: begin
				q			<=			16'hFFFF;
		end
		32'h0000F938: begin
				q			<=			16'hD7D0;
		end
		32'h0000F93A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F93C: begin
				q			<=			16'hD784;
		end
		32'h0000F93E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F940: begin
				q			<=			16'hD784;
		end
		32'h0000F942: begin
				q			<=			16'hFFFF;
		end
		32'h0000F944: begin
				q			<=			16'hDA44;
		end
		32'h0000F946: begin
				q			<=			16'hFFFF;
		end
		32'h0000F948: begin
				q			<=			16'hD7D0;
		end
		32'h0000F94A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F94C: begin
				q			<=			16'hD784;
		end
		32'h0000F94E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F950: begin
				q			<=			16'hDA44;
		end
		32'h0000F952: begin
				q			<=			16'hFFFF;
		end
		32'h0000F954: begin
				q			<=			16'hD784;
		end
		32'h0000F956: begin
				q			<=			16'hFFFF;
		end
		32'h0000F958: begin
				q			<=			16'hD7D0;
		end
		32'h0000F95A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F95C: begin
				q			<=			16'hD780;
		end
		32'h0000F95E: begin
				q			<=			16'hFFFF;
		end
		32'h0000F960: begin
				q			<=			16'hD780;
		end
		32'h0000F962: begin
				q			<=			16'hFFFF;
		end
		32'h0000F964: begin
				q			<=			16'hD780;
		end
		32'h0000F966: begin
				q			<=			16'hFFFF;
		end
		32'h0000F968: begin
				q			<=			16'hDA44;
		end
		32'h0000F96A: begin
				q			<=			16'hFFFF;
		end
		32'h0000F96C: begin
				q			<=			16'h0100;
		end
		32'h0000F96E: begin
				q			<=			16'h0202;
		end
		32'h0000F970: begin
				q			<=			16'h0303;
		end
		32'h0000F972: begin
				q			<=			16'h0303;
		end
		32'h0000F974: begin
				q			<=			16'h0404;
		end
		32'h0000F976: begin
				q			<=			16'h0404;
		end
		32'h0000F978: begin
				q			<=			16'h0404;
		end
		32'h0000F97A: begin
				q			<=			16'h0404;
		end
		32'h0000F97C: begin
				q			<=			16'h0505;
		end
		32'h0000F97E: begin
				q			<=			16'h0505;
		end
		32'h0000F980: begin
				q			<=			16'h0505;
		end
		32'h0000F982: begin
				q			<=			16'h0505;
		end
		32'h0000F984: begin
				q			<=			16'h0505;
		end
		32'h0000F986: begin
				q			<=			16'h0505;
		end
		32'h0000F988: begin
				q			<=			16'h0505;
		end
		32'h0000F98A: begin
				q			<=			16'h0505;
		end
		32'h0000F98C: begin
				q			<=			16'h0606;
		end
		32'h0000F98E: begin
				q			<=			16'h0606;
		end
		32'h0000F990: begin
				q			<=			16'h0606;
		end
		32'h0000F992: begin
				q			<=			16'h0606;
		end
		32'h0000F994: begin
				q			<=			16'h0606;
		end
		32'h0000F996: begin
				q			<=			16'h0606;
		end
		32'h0000F998: begin
				q			<=			16'h0606;
		end
		32'h0000F99A: begin
				q			<=			16'h0606;
		end
		32'h0000F99C: begin
				q			<=			16'h0606;
		end
		32'h0000F99E: begin
				q			<=			16'h0606;
		end
		32'h0000F9A0: begin
				q			<=			16'h0606;
		end
		32'h0000F9A2: begin
				q			<=			16'h0606;
		end
		32'h0000F9A4: begin
				q			<=			16'h0606;
		end
		32'h0000F9A6: begin
				q			<=			16'h0606;
		end
		32'h0000F9A8: begin
				q			<=			16'h0606;
		end
		32'h0000F9AA: begin
				q			<=			16'h0606;
		end
		32'h0000F9AC: begin
				q			<=			16'h0707;
		end
		32'h0000F9AE: begin
				q			<=			16'h0707;
		end
		32'h0000F9B0: begin
				q			<=			16'h0707;
		end
		32'h0000F9B2: begin
				q			<=			16'h0707;
		end
		32'h0000F9B4: begin
				q			<=			16'h0707;
		end
		32'h0000F9B6: begin
				q			<=			16'h0707;
		end
		32'h0000F9B8: begin
				q			<=			16'h0707;
		end
		32'h0000F9BA: begin
				q			<=			16'h0707;
		end
		32'h0000F9BC: begin
				q			<=			16'h0707;
		end
		32'h0000F9BE: begin
				q			<=			16'h0707;
		end
		32'h0000F9C0: begin
				q			<=			16'h0707;
		end
		32'h0000F9C2: begin
				q			<=			16'h0707;
		end
		32'h0000F9C4: begin
				q			<=			16'h0707;
		end
		32'h0000F9C6: begin
				q			<=			16'h0707;
		end
		32'h0000F9C8: begin
				q			<=			16'h0707;
		end
		32'h0000F9CA: begin
				q			<=			16'h0707;
		end
		32'h0000F9CC: begin
				q			<=			16'h0707;
		end
		32'h0000F9CE: begin
				q			<=			16'h0707;
		end
		32'h0000F9D0: begin
				q			<=			16'h0707;
		end
		32'h0000F9D2: begin
				q			<=			16'h0707;
		end
		32'h0000F9D4: begin
				q			<=			16'h0707;
		end
		32'h0000F9D6: begin
				q			<=			16'h0707;
		end
		32'h0000F9D8: begin
				q			<=			16'h0707;
		end
		32'h0000F9DA: begin
				q			<=			16'h0707;
		end
		32'h0000F9DC: begin
				q			<=			16'h0707;
		end
		32'h0000F9DE: begin
				q			<=			16'h0707;
		end
		32'h0000F9E0: begin
				q			<=			16'h0707;
		end
		32'h0000F9E2: begin
				q			<=			16'h0707;
		end
		32'h0000F9E4: begin
				q			<=			16'h0707;
		end
		32'h0000F9E6: begin
				q			<=			16'h0707;
		end
		32'h0000F9E8: begin
				q			<=			16'h0707;
		end
		32'h0000F9EA: begin
				q			<=			16'h0707;
		end
		32'h0000F9EC: begin
				q			<=			16'h0808;
		end
		32'h0000F9EE: begin
				q			<=			16'h0808;
		end
		32'h0000F9F0: begin
				q			<=			16'h0808;
		end
		32'h0000F9F2: begin
				q			<=			16'h0808;
		end
		32'h0000F9F4: begin
				q			<=			16'h0808;
		end
		32'h0000F9F6: begin
				q			<=			16'h0808;
		end
		32'h0000F9F8: begin
				q			<=			16'h0808;
		end
		32'h0000F9FA: begin
				q			<=			16'h0808;
		end
		32'h0000F9FC: begin
				q			<=			16'h0808;
		end
		32'h0000F9FE: begin
				q			<=			16'h0808;
		end
		32'h0000FA00: begin
				q			<=			16'h0808;
		end
		32'h0000FA02: begin
				q			<=			16'h0808;
		end
		32'h0000FA04: begin
				q			<=			16'h0808;
		end
		32'h0000FA06: begin
				q			<=			16'h0808;
		end
		32'h0000FA08: begin
				q			<=			16'h0808;
		end
		32'h0000FA0A: begin
				q			<=			16'h0808;
		end
		32'h0000FA0C: begin
				q			<=			16'h0808;
		end
		32'h0000FA0E: begin
				q			<=			16'h0808;
		end
		32'h0000FA10: begin
				q			<=			16'h0808;
		end
		32'h0000FA12: begin
				q			<=			16'h0808;
		end
		32'h0000FA14: begin
				q			<=			16'h0808;
		end
		32'h0000FA16: begin
				q			<=			16'h0808;
		end
		32'h0000FA18: begin
				q			<=			16'h0808;
		end
		32'h0000FA1A: begin
				q			<=			16'h0808;
		end
		32'h0000FA1C: begin
				q			<=			16'h0808;
		end
		32'h0000FA1E: begin
				q			<=			16'h0808;
		end
		32'h0000FA20: begin
				q			<=			16'h0808;
		end
		32'h0000FA22: begin
				q			<=			16'h0808;
		end
		32'h0000FA24: begin
				q			<=			16'h0808;
		end
		32'h0000FA26: begin
				q			<=			16'h0808;
		end
		32'h0000FA28: begin
				q			<=			16'h0808;
		end
		32'h0000FA2A: begin
				q			<=			16'h0808;
		end
		32'h0000FA2C: begin
				q			<=			16'h0808;
		end
		32'h0000FA2E: begin
				q			<=			16'h0808;
		end
		32'h0000FA30: begin
				q			<=			16'h0808;
		end
		32'h0000FA32: begin
				q			<=			16'h0808;
		end
		32'h0000FA34: begin
				q			<=			16'h0808;
		end
		32'h0000FA36: begin
				q			<=			16'h0808;
		end
		32'h0000FA38: begin
				q			<=			16'h0808;
		end
		32'h0000FA3A: begin
				q			<=			16'h0808;
		end
		32'h0000FA3C: begin
				q			<=			16'h0808;
		end
		32'h0000FA3E: begin
				q			<=			16'h0808;
		end
		32'h0000FA40: begin
				q			<=			16'h0808;
		end
		32'h0000FA42: begin
				q			<=			16'h0808;
		end
		32'h0000FA44: begin
				q			<=			16'h0808;
		end
		32'h0000FA46: begin
				q			<=			16'h0808;
		end
		32'h0000FA48: begin
				q			<=			16'h0808;
		end
		32'h0000FA4A: begin
				q			<=			16'h0808;
		end
		32'h0000FA4C: begin
				q			<=			16'h0808;
		end
		32'h0000FA4E: begin
				q			<=			16'h0808;
		end
		32'h0000FA50: begin
				q			<=			16'h0808;
		end
		32'h0000FA52: begin
				q			<=			16'h0808;
		end
		32'h0000FA54: begin
				q			<=			16'h0808;
		end
		32'h0000FA56: begin
				q			<=			16'h0808;
		end
		32'h0000FA58: begin
				q			<=			16'h0808;
		end
		32'h0000FA5A: begin
				q			<=			16'h0808;
		end
		32'h0000FA5C: begin
				q			<=			16'h0808;
		end
		32'h0000FA5E: begin
				q			<=			16'h0808;
		end
		32'h0000FA60: begin
				q			<=			16'h0808;
		end
		32'h0000FA62: begin
				q			<=			16'h0808;
		end
		32'h0000FA64: begin
				q			<=			16'h0808;
		end
		32'h0000FA66: begin
				q			<=			16'h0808;
		end
		32'h0000FA68: begin
				q			<=			16'h0808;
		end
		32'h0000FA6A: begin
				q			<=			16'h0808;
		end
		32'h0000FA6C: begin
				q			<=			16'h435B;
		end
		32'h0000FA6E: begin
				q			<=			16'h4E4F;
		end
		32'h0000FA70: begin
				q			<=			16'h4F53;
		end
		32'h0000FA72: begin
				q			<=			16'h454C;
		end
		32'h0000FA74: begin
				q			<=			16'h4320;
		end
		32'h0000FA76: begin
				q			<=			16'h4D4F;
		end
		32'h0000FA78: begin
				q			<=			16'h414D;
		end
		32'h0000FA7A: begin
				q			<=			16'h444E;
		end
		32'h0000FA7C: begin
				q			<=			16'h4C20;
		end
		32'h0000FA7E: begin
				q			<=			16'h5349;
		end
		32'h0000FA80: begin
				q			<=			16'h5D54;
		end
		32'h0000FA82: begin
				q			<=			16'h0000;
		end
		32'h0000FA84: begin
				q			<=			16'h4C43;
		end
		32'h0000FA86: begin
				q			<=			16'h2053;
		end
		32'h0000FA88: begin
				q			<=			16'h2020;
		end
		32'h0000FA8A: begin
				q			<=			16'h2020;
		end
		32'h0000FA8C: begin
				q			<=			16'h2020;
		end
		32'h0000FA8E: begin
				q			<=			16'h2020;
		end
		32'h0000FA90: begin
				q			<=			16'h2020;
		end
		32'h0000FA92: begin
				q			<=			16'h4320;
		end
		32'h0000FA94: begin
				q			<=			16'h454C;
		end
		32'h0000FA96: begin
				q			<=			16'h5241;
		end
		32'h0000FA98: begin
				q			<=			16'h5320;
		end
		32'h0000FA9A: begin
				q			<=			16'h5243;
		end
		32'h0000FA9C: begin
				q			<=			16'h4545;
		end
		32'h0000FA9E: begin
				q			<=			16'h204E;
		end
		32'h0000FAA0: begin
				q			<=			16'h4554;
		end
		32'h0000FAA2: begin
				q			<=			16'h5458;
		end
		32'h0000FAA4: begin
				q			<=			16'h0000;
		end
		32'h0000FAA6: begin
				q			<=			16'h0000;
		end
		32'h0000FAA8: begin
				q			<=			16'h4443;
		end
		32'h0000FAAA: begin
				q			<=			16'h7820;
		end
		32'h0000FAAC: begin
				q			<=			16'h2020;
		end
		32'h0000FAAE: begin
				q			<=			16'h2020;
		end
		32'h0000FAB0: begin
				q			<=			16'h2020;
		end
		32'h0000FAB2: begin
				q			<=			16'h2020;
		end
		32'h0000FAB4: begin
				q			<=			16'h2020;
		end
		32'h0000FAB6: begin
				q			<=			16'h4320;
		end
		32'h0000FAB8: begin
				q			<=			16'h4148;
		end
		32'h0000FABA: begin
				q			<=			16'h474E;
		end
		32'h0000FABC: begin
				q			<=			16'h2045;
		end
		32'h0000FABE: begin
				q			<=			16'h4944;
		end
		32'h0000FAC0: begin
				q			<=			16'h4552;
		end
		32'h0000FAC2: begin
				q			<=			16'h5443;
		end
		32'h0000FAC4: begin
				q			<=			16'h524F;
		end
		32'h0000FAC6: begin
				q			<=			16'h0059;
		end
		32'h0000FAC8: begin
				q			<=			16'h4944;
		end
		32'h0000FACA: begin
				q			<=			16'h2052;
		end
		32'h0000FACC: begin
				q			<=			16'h2020;
		end
		32'h0000FACE: begin
				q			<=			16'h2020;
		end
		32'h0000FAD0: begin
				q			<=			16'h2020;
		end
		32'h0000FAD2: begin
				q			<=			16'h2020;
		end
		32'h0000FAD4: begin
				q			<=			16'h2020;
		end
		32'h0000FAD6: begin
				q			<=			16'h4C20;
		end
		32'h0000FAD8: begin
				q			<=			16'h5349;
		end
		32'h0000FADA: begin
				q			<=			16'h2054;
		end
		32'h0000FADC: begin
				q			<=			16'h4944;
		end
		32'h0000FADE: begin
				q			<=			16'h4552;
		end
		32'h0000FAE0: begin
				q			<=			16'h5443;
		end
		32'h0000FAE2: begin
				q			<=			16'h524F;
		end
		32'h0000FAE4: begin
				q			<=			16'h0059;
		end
		32'h0000FAE6: begin
				q			<=			16'h0000;
		end
		32'h0000FAE8: begin
				q			<=			16'h5753;
		end
		32'h0000FAEA: begin
				q			<=			16'h5041;
		end
		32'h0000FAEC: begin
				q			<=			16'h464F;
		end
		32'h0000FAEE: begin
				q			<=			16'h2046;
		end
		32'h0000FAF0: begin
				q			<=			16'h2020;
		end
		32'h0000FAF2: begin
				q			<=			16'h2020;
		end
		32'h0000FAF4: begin
				q			<=			16'h2020;
		end
		32'h0000FAF6: begin
				q			<=			16'h4120;
		end
		32'h0000FAF8: begin
				q			<=			16'h5455;
		end
		32'h0000FAFA: begin
				q			<=			16'h204F;
		end
		32'h0000FAFC: begin
				q			<=			16'h4F44;
		end
		32'h0000FAFE: begin
				q			<=			16'h4255;
		end
		32'h0000FB00: begin
				q			<=			16'h454C;
		end
		32'h0000FB02: begin
				q			<=			16'h4220;
		end
		32'h0000FB04: begin
				q			<=			16'h4655;
		end
		32'h0000FB06: begin
				q			<=			16'h4546;
		end
		32'h0000FB08: begin
				q			<=			16'h2052;
		end
		32'h0000FB0A: begin
				q			<=			16'h5753;
		end
		32'h0000FB0C: begin
				q			<=			16'h5041;
		end
		32'h0000FB0E: begin
				q			<=			16'h4F20;
		end
		32'h0000FB10: begin
				q			<=			16'h4646;
		end
		32'h0000FB12: begin
				q			<=			16'h0000;
		end
		32'h0000FB14: begin
				q			<=			16'h5753;
		end
		32'h0000FB16: begin
				q			<=			16'h5041;
		end
		32'h0000FB18: begin
				q			<=			16'h4E4F;
		end
		32'h0000FB1A: begin
				q			<=			16'h2020;
		end
		32'h0000FB1C: begin
				q			<=			16'h2020;
		end
		32'h0000FB1E: begin
				q			<=			16'h2020;
		end
		32'h0000FB20: begin
				q			<=			16'h2020;
		end
		32'h0000FB22: begin
				q			<=			16'h4120;
		end
		32'h0000FB24: begin
				q			<=			16'h5455;
		end
		32'h0000FB26: begin
				q			<=			16'h204F;
		end
		32'h0000FB28: begin
				q			<=			16'h4F44;
		end
		32'h0000FB2A: begin
				q			<=			16'h4255;
		end
		32'h0000FB2C: begin
				q			<=			16'h454C;
		end
		32'h0000FB2E: begin
				q			<=			16'h4220;
		end
		32'h0000FB30: begin
				q			<=			16'h4655;
		end
		32'h0000FB32: begin
				q			<=			16'h4546;
		end
		32'h0000FB34: begin
				q			<=			16'h2052;
		end
		32'h0000FB36: begin
				q			<=			16'h5753;
		end
		32'h0000FB38: begin
				q			<=			16'h5041;
		end
		32'h0000FB3A: begin
				q			<=			16'h4F20;
		end
		32'h0000FB3C: begin
				q			<=			16'h004E;
		end
		32'h0000FB3E: begin
				q			<=			16'h0000;
		end
		32'h0000FB40: begin
				q			<=			16'h5753;
		end
		32'h0000FB42: begin
				q			<=			16'h5041;
		end
		32'h0000FB44: begin
				q			<=			16'h4F4E;
		end
		32'h0000FB46: begin
				q			<=			16'h2057;
		end
		32'h0000FB48: begin
				q			<=			16'h2020;
		end
		32'h0000FB4A: begin
				q			<=			16'h2020;
		end
		32'h0000FB4C: begin
				q			<=			16'h2020;
		end
		32'h0000FB4E: begin
				q			<=			16'h5320;
		end
		32'h0000FB50: begin
				q			<=			16'h4157;
		end
		32'h0000FB52: begin
				q			<=			16'h2050;
		end
		32'h0000FB54: begin
				q			<=			16'h4F44;
		end
		32'h0000FB56: begin
				q			<=			16'h4255;
		end
		32'h0000FB58: begin
				q			<=			16'h454C;
		end
		32'h0000FB5A: begin
				q			<=			16'h4220;
		end
		32'h0000FB5C: begin
				q			<=			16'h4655;
		end
		32'h0000FB5E: begin
				q			<=			16'h4546;
		end
		32'h0000FB60: begin
				q			<=			16'h5352;
		end
		32'h0000FB62: begin
				q			<=			16'h4E20;
		end
		32'h0000FB64: begin
				q			<=			16'h574F;
		end
		32'h0000FB66: begin
				q			<=			16'h0000;
		end
		32'h0000FB68: begin
				q			<=			16'h4C42;
		end
		32'h0000FB6A: begin
				q			<=			16'h4341;
		end
		32'h0000FB6C: begin
				q			<=			16'h424B;
		end
		32'h0000FB6E: begin
				q			<=			16'h4655;
		end
		32'h0000FB70: begin
				q			<=			16'h2020;
		end
		32'h0000FB72: begin
				q			<=			16'h2020;
		end
		32'h0000FB74: begin
				q			<=			16'h2020;
		end
		32'h0000FB76: begin
				q			<=			16'h4220;
		end
		32'h0000FB78: begin
				q			<=			16'h414C;
		end
		32'h0000FB7A: begin
				q			<=			16'h4B43;
		end
		32'h0000FB7C: begin
				q			<=			16'h4320;
		end
		32'h0000FB7E: begin
				q			<=			16'h5255;
		end
		32'h0000FB80: begin
				q			<=			16'h4552;
		end
		32'h0000FB82: begin
				q			<=			16'h544E;
		end
		32'h0000FB84: begin
				q			<=			16'h4220;
		end
		32'h0000FB86: begin
				q			<=			16'h4655;
		end
		32'h0000FB88: begin
				q			<=			16'h4546;
		end
		32'h0000FB8A: begin
				q			<=			16'h0052;
		end
		32'h0000FB8C: begin
				q			<=			16'h4857;
		end
		32'h0000FB8E: begin
				q			<=			16'h5449;
		end
		32'h0000FB90: begin
				q			<=			16'h4245;
		end
		32'h0000FB92: begin
				q			<=			16'h4655;
		end
		32'h0000FB94: begin
				q			<=			16'h2020;
		end
		32'h0000FB96: begin
				q			<=			16'h2020;
		end
		32'h0000FB98: begin
				q			<=			16'h2020;
		end
		32'h0000FB9A: begin
				q			<=			16'h5720;
		end
		32'h0000FB9C: begin
				q			<=			16'h4948;
		end
		32'h0000FB9E: begin
				q			<=			16'h4554;
		end
		32'h0000FBA0: begin
				q			<=			16'h4320;
		end
		32'h0000FBA2: begin
				q			<=			16'h5255;
		end
		32'h0000FBA4: begin
				q			<=			16'h4552;
		end
		32'h0000FBA6: begin
				q			<=			16'h544E;
		end
		32'h0000FBA8: begin
				q			<=			16'h4220;
		end
		32'h0000FBAA: begin
				q			<=			16'h4655;
		end
		32'h0000FBAC: begin
				q			<=			16'h4546;
		end
		32'h0000FBAE: begin
				q			<=			16'h0052;
		end
		32'h0000FBB0: begin
				q			<=			16'h4548;
		end
		32'h0000FBB2: begin
				q			<=			16'h504C;
		end
		32'h0000FBB4: begin
				q			<=			16'h0000;
		end
		32'h0000FBB6: begin
				q			<=			16'h0000;
		end
		32'h0000FBB8: begin
				q			<=			16'h4C43;
		end
		32'h0000FBBA: begin
				q			<=			16'h0053;
		end
		32'h0000FBBC: begin
				q			<=			16'h4944;
		end
		32'h0000FBBE: begin
				q			<=			16'h0052;
		end
		32'h0000FBC0: begin
				q			<=			16'h4443;
		end
		32'h0000FBC2: begin
				q			<=			16'h0020;
		end
		32'h0000FBC4: begin
				q			<=			16'h504F;
		end
		32'h0000FBC6: begin
				q			<=			16'h4E45;
		end
		32'h0000FBC8: begin
				q			<=			16'h4420;
		end
		32'h0000FBCA: begin
				q			<=			16'h5249;
		end
		32'h0000FBCC: begin
				q			<=			16'h4345;
		end
		32'h0000FBCE: begin
				q			<=			16'h4F54;
		end
		32'h0000FBD0: begin
				q			<=			16'h5952;
		end
		32'h0000FBD2: begin
				q			<=			16'h4520;
		end
		32'h0000FBD4: begin
				q			<=			16'h5252;
		end
		32'h0000FBD6: begin
				q			<=			16'h524F;
		end
		32'h0000FBD8: begin
				q			<=			16'h0021;
		end
		32'h0000FBDA: begin
				q			<=			16'h0000;
		end
		32'h0000FBDC: begin
				q			<=			16'h504F;
		end
		32'h0000FBDE: begin
				q			<=			16'h4E45;
		end
		32'h0000FBE0: begin
				q			<=			16'h4420;
		end
		32'h0000FBE2: begin
				q			<=			16'h5249;
		end
		32'h0000FBE4: begin
				q			<=			16'h4345;
		end
		32'h0000FBE6: begin
				q			<=			16'h4F54;
		end
		32'h0000FBE8: begin
				q			<=			16'h5952;
		end
		32'h0000FBEA: begin
				q			<=			16'h5320;
		end
		32'h0000FBEC: begin
				q			<=			16'h4355;
		end
		32'h0000FBEE: begin
				q			<=			16'h4543;
		end
		32'h0000FBF0: begin
				q			<=			16'h5353;
		end
		32'h0000FBF2: begin
				q			<=			16'h0000;
		end
		32'h0000FBF4: begin
				q			<=			16'h4C42;
		end
		32'h0000FBF6: begin
				q			<=			16'h4341;
		end
		32'h0000FBF8: begin
				q			<=			16'h424B;
		end
		32'h0000FBFA: begin
				q			<=			16'h4655;
		end
		32'h0000FBFC: begin
				q			<=			16'h0000;
		end
		32'h0000FBFE: begin
				q			<=			16'h0000;
		end
		32'h0000FC00: begin
				q			<=			16'h5542;
		end
		32'h0000FC02: begin
				q			<=			16'h4646;
		end
		32'h0000FC04: begin
				q			<=			16'h5245;
		end
		32'h0000FC06: begin
				q			<=			16'h4220;
		end
		32'h0000FC08: begin
				q			<=			16'h414C;
		end
		32'h0000FC0A: begin
				q			<=			16'h4B43;
		end
		32'h0000FC0C: begin
				q			<=			16'h4445;
		end
		32'h0000FC0E: begin
				q			<=			16'h0000;
		end
		32'h0000FC10: begin
				q			<=			16'h4857;
		end
		32'h0000FC12: begin
				q			<=			16'h5449;
		end
		32'h0000FC14: begin
				q			<=			16'h4245;
		end
		32'h0000FC16: begin
				q			<=			16'h4655;
		end
		32'h0000FC18: begin
				q			<=			16'h0000;
		end
		32'h0000FC1A: begin
				q			<=			16'h0000;
		end
		32'h0000FC1C: begin
				q			<=			16'h5542;
		end
		32'h0000FC1E: begin
				q			<=			16'h4646;
		end
		32'h0000FC20: begin
				q			<=			16'h5245;
		end
		32'h0000FC22: begin
				q			<=			16'h5720;
		end
		32'h0000FC24: begin
				q			<=			16'h4948;
		end
		32'h0000FC26: begin
				q			<=			16'h4554;
		end
		32'h0000FC28: begin
				q			<=			16'h0044;
		end
		32'h0000FC2A: begin
				q			<=			16'h0000;
		end
		32'h0000FC2C: begin
				q			<=			16'h5753;
		end
		32'h0000FC2E: begin
				q			<=			16'h5041;
		end
		32'h0000FC30: begin
				q			<=			16'h464F;
		end
		32'h0000FC32: begin
				q			<=			16'h0046;
		end
		32'h0000FC34: begin
				q			<=			16'h5541;
		end
		32'h0000FC36: begin
				q			<=			16'h4F54;
		end
		32'h0000FC38: begin
				q			<=			16'h5320;
		end
		32'h0000FC3A: begin
				q			<=			16'h4157;
		end
		32'h0000FC3C: begin
				q			<=			16'h2050;
		end
		32'h0000FC3E: begin
				q			<=			16'h464F;
		end
		32'h0000FC40: begin
				q			<=			16'h0046;
		end
		32'h0000FC42: begin
				q			<=			16'h0000;
		end
		32'h0000FC44: begin
				q			<=			16'h5753;
		end
		32'h0000FC46: begin
				q			<=			16'h5041;
		end
		32'h0000FC48: begin
				q			<=			16'h4E4F;
		end
		32'h0000FC4A: begin
				q			<=			16'h0000;
		end
		32'h0000FC4C: begin
				q			<=			16'h5753;
		end
		32'h0000FC4E: begin
				q			<=			16'h5041;
		end
		32'h0000FC50: begin
				q			<=			16'h4F4E;
		end
		32'h0000FC52: begin
				q			<=			16'h0057;
		end
		32'h0000FC54: begin
				q			<=			16'h5753;
		end
		32'h0000FC56: begin
				q			<=			16'h5041;
		end
		32'h0000FC58: begin
				q			<=			16'h4550;
		end
		32'h0000FC5A: begin
				q			<=			16'h2044;
		end
		32'h0000FC5C: begin
				q			<=			16'h4F54;
		end
		32'h0000FC5E: begin
				q			<=			16'h4220;
		end
		32'h0000FC60: begin
				q			<=			16'h4220;
		end
		32'h0000FC62: begin
				q			<=			16'h4655;
		end
		32'h0000FC64: begin
				q			<=			16'h4546;
		end
		32'h0000FC66: begin
				q			<=			16'h0052;
		end
		32'h0000FC68: begin
				q			<=			16'h5753;
		end
		32'h0000FC6A: begin
				q			<=			16'h5041;
		end
		32'h0000FC6C: begin
				q			<=			16'h4550;
		end
		32'h0000FC6E: begin
				q			<=			16'h2044;
		end
		32'h0000FC70: begin
				q			<=			16'h4F54;
		end
		32'h0000FC72: begin
				q			<=			16'h4120;
		end
		32'h0000FC74: begin
				q			<=			16'h4220;
		end
		32'h0000FC76: begin
				q			<=			16'h4655;
		end
		32'h0000FC78: begin
				q			<=			16'h4546;
		end
		32'h0000FC7A: begin
				q			<=			16'h0052;
		end
		32'h0000FC7C: begin
				q			<=			16'h5453;
		end
		32'h0000FC7E: begin
				q			<=			16'h5441;
		end
		32'h0000FC80: begin
				q			<=			16'h5355;
		end
		32'h0000FC82: begin
				q			<=			16'h0000;
		end
		32'h0000FC84: begin
				q			<=			16'h5453;
		end
		32'h0000FC86: begin
				q			<=			16'h5441;
		end
		32'h0000FC88: begin
				q			<=			16'h5355;
		end
		32'h0000FC8A: begin
				q			<=			16'h2D20;
		end
		32'h0000FC8C: begin
				q			<=			16'h0020;
		end
		32'h0000FC8E: begin
				q			<=			16'h0000;
		end
		32'h0000FC90: begin
				q			<=			16'h535B;
		end
		32'h0000FC92: begin
				q			<=			16'h5359;
		end
		32'h0000FC94: begin
				q			<=			16'h4554;
		end
		32'h0000FC96: begin
				q			<=			16'h5D4D;
		end
		32'h0000FC98: begin
				q			<=			16'h0020;
		end
		32'h0000FC9A: begin
				q			<=			16'h0000;
		end
		32'h0000FC9C: begin
				q			<=			16'h7325;
		end
		32'h0000FC9E: begin
				q			<=			16'h2520;
		end
		32'h0000FCA0: begin
				q			<=			16'h0073;
		end
		32'h0000FCA2: begin
				q			<=			16'h0000;
		end
		32'h0000FCA4: begin
				q			<=			16'h7325;
		end
		32'h0000FCA6: begin
				q			<=			16'h7325;
		end
		32'h0000FCA8: begin
				q			<=			16'h7325;
		end
		32'h0000FCAA: begin
				q			<=			16'h7325;
		end
		32'h0000FCAC: begin
				q			<=			16'h7325;
		end
		32'h0000FCAE: begin
				q			<=			16'h7325;
		end
		32'h0000FCB0: begin
				q			<=			16'h7325;
		end
		32'h0000FCB2: begin
				q			<=			16'h7325;
		end
		32'h0000FCB4: begin
				q			<=			16'h0000;
		end
		32'h0000FCB6: begin
				q			<=			16'h0000;
		end
		32'h0000FCB8: begin
				q			<=			16'h7325;
		end
		32'h0000FCBA: begin
				q			<=			16'h7325;
		end
		32'h0000FCBC: begin
				q			<=			16'h7325;
		end
		32'h0000FCBE: begin
				q			<=			16'h7325;
		end
		32'h0000FCC0: begin
				q			<=			16'h7325;
		end
		32'h0000FCC2: begin
				q			<=			16'h7325;
		end
		32'h0000FCC4: begin
				q			<=			16'h7325;
		end
		32'h0000FCC6: begin
				q			<=			16'h7325;
		end
		32'h0000FCC8: begin
				q			<=			16'h7325;
		end
		32'h0000FCCA: begin
				q			<=			16'h0000;
		end
		32'h0000FCCC: begin
				q			<=			16'h7830;
		end
		32'h0000FCCE: begin
				q			<=			16'h2530;
		end
		32'h0000FCD0: begin
				q			<=			16'h3830;
		end
		32'h0000FCD2: begin
				q			<=			16'h0078;
		end
		32'h0000FCD4: begin
				q			<=			16'h1324;
		end
		32'h0000FCD6: begin
				q			<=			16'h0000;
		end
		32'h0000FCD8: begin
				q			<=			16'h1340;
		end
		32'h0000FCDA: begin
				q			<=			16'h0000;
		end
		32'h0000FCDC: begin
				q			<=			16'h1354;
		end
		32'h0000FCDE: begin
				q			<=			16'h0000;
		end
		32'h0000FCE0: begin
				q			<=			16'h1368;
		end
		32'h0000FCE2: begin
				q			<=			16'h0000;
		end
		32'h0000FCE4: begin
				q			<=			16'h137C;
		end
		32'h0000FCE6: begin
				q			<=			16'h0000;
		end
		32'h0000FCE8: begin
				q			<=			16'h465B;
		end
		32'h0000FCEA: begin
				q			<=			16'h6961;
		end
		32'h0000FCEC: begin
				q			<=			16'h206C;
		end
		32'h0000FCEE: begin
				q			<=			16'h6372;
		end
		32'h0000FCF0: begin
				q			<=			16'h253D;
		end
		32'h0000FCF2: begin
				q			<=			16'h5D75;
		end
		32'h0000FCF4: begin
				q			<=			16'h0000;
		end
		32'h0000FCF6: begin
				q			<=			16'h0000;
		end
		32'h0000FCF8: begin
				q			<=			16'h4F4E;
		end
		32'h0000FCFA: begin
				q			<=			16'h4520;
		end
		32'h0000FCFC: begin
				q			<=			16'h5252;
		end
		32'h0000FCFE: begin
				q			<=			16'h524F;
		end
		32'h0000FD00: begin
				q			<=			16'h0000;
		end
		32'h0000FD02: begin
				q			<=			16'h0000;
		end
		32'h0000FD04: begin
				q			<=			16'h4946;
		end
		32'h0000FD06: begin
				q			<=			16'h454C;
		end
		32'h0000FD08: begin
				q			<=			16'h5320;
		end
		32'h0000FD0A: begin
				q			<=			16'h5359;
		end
		32'h0000FD0C: begin
				q			<=			16'h4554;
		end
		32'h0000FD0E: begin
				q			<=			16'h204D;
		end
		32'h0000FD10: begin
				q			<=			16'h5245;
		end
		32'h0000FD12: begin
				q			<=			16'h4F52;
		end
		32'h0000FD14: begin
				q			<=			16'h0052;
		end
		32'h0000FD16: begin
				q			<=			16'h0000;
		end
		32'h0000FD18: begin
				q			<=			16'h4946;
		end
		32'h0000FD1A: begin
				q			<=			16'h454C;
		end
		32'h0000FD1C: begin
				q			<=			16'h4920;
		end
		32'h0000FD1E: begin
				q			<=			16'h204F;
		end
		32'h0000FD20: begin
				q			<=			16'h5245;
		end
		32'h0000FD22: begin
				q			<=			16'h4F52;
		end
		32'h0000FD24: begin
				q			<=			16'h0052;
		end
		32'h0000FD26: begin
				q			<=			16'h0000;
		end
		32'h0000FD28: begin
				q			<=			16'h5247;
		end
		32'h0000FD2A: begin
				q			<=			16'h5041;
		end
		32'h0000FD2C: begin
				q			<=			16'h4948;
		end
		32'h0000FD2E: begin
				q			<=			16'h5343;
		end
		32'h0000FD30: begin
				q			<=			16'h4920;
		end
		32'h0000FD32: begin
				q			<=			16'h204F;
		end
		32'h0000FD34: begin
				q			<=			16'h5245;
		end
		32'h0000FD36: begin
				q			<=			16'h4F52;
		end
		32'h0000FD38: begin
				q			<=			16'h0052;
		end
		32'h0000FD3A: begin
				q			<=			16'h0000;
		end
		32'h0000FD3C: begin
				q			<=			16'h454D;
		end
		32'h0000FD3E: begin
				q			<=			16'h4F4D;
		end
		32'h0000FD40: begin
				q			<=			16'h5952;
		end
		32'h0000FD42: begin
				q			<=			16'h4520;
		end
		32'h0000FD44: begin
				q			<=			16'h5252;
		end
		32'h0000FD46: begin
				q			<=			16'h524F;
		end
		32'h0000FD48: begin
				q			<=			16'h0000;
		end
		32'h0000FD4A: begin
				q			<=			16'h0000;
		end
		32'h0000FD4C: begin
				q			<=			16'h4E55;
		end
		32'h0000FD4E: begin
				q			<=			16'h4E4B;
		end
		32'h0000FD50: begin
				q			<=			16'h574F;
		end
		32'h0000FD52: begin
				q			<=			16'h204E;
		end
		32'h0000FD54: begin
				q			<=			16'h5245;
		end
		32'h0000FD56: begin
				q			<=			16'h4F52;
		end
		32'h0000FD58: begin
				q			<=			16'h0052;
		end
		32'h0000FD5A: begin
				q			<=			16'h0000;
		end
		32'h0000FD5C: begin
				q			<=			16'h443C;
		end
		32'h0000FD5E: begin
				q			<=			16'h5249;
		end
		32'h0000FD60: begin
				q			<=			16'h203E;
		end
		32'h0000FD62: begin
				q			<=			16'h7325;
		end
		32'h0000FD64: begin
				q			<=			16'h0000;
		end
		32'h0000FD66: begin
				q			<=			16'h0000;
		end
		32'h0000FD68: begin
				q			<=			16'h2020;
		end
		32'h0000FD6A: begin
				q			<=			16'h2020;
		end
		32'h0000FD6C: begin
				q			<=			16'h2020;
		end
		32'h0000FD6E: begin
				q			<=			16'h7325;
		end
		32'h0000FD70: begin
				q			<=			16'h0000;
		end
		32'h0000FD72: begin
				q			<=			16'h0000;
		end
		32'h0000FD74: begin
				q			<=			16'h4E49;
		end
		32'h0000FD76: begin
				q			<=			16'h0046;
		end
		32'h0000FD78: begin
				q			<=			16'h6E69;
		end
		32'h0000FD7A: begin
				q			<=			16'h0066;
		end
		32'h0000FD7C: begin
				q			<=			16'h414E;
		end
		32'h0000FD7E: begin
				q			<=			16'h004E;
		end
		32'h0000FD80: begin
				q			<=			16'h616E;
		end
		32'h0000FD82: begin
				q			<=			16'h006E;
		end
		32'h0000FD84: begin
				q			<=			16'h3130;
		end
		32'h0000FD86: begin
				q			<=			16'h3332;
		end
		32'h0000FD88: begin
				q			<=			16'h3534;
		end
		32'h0000FD8A: begin
				q			<=			16'h3736;
		end
		32'h0000FD8C: begin
				q			<=			16'h3938;
		end
		32'h0000FD8E: begin
				q			<=			16'h6261;
		end
		32'h0000FD90: begin
				q			<=			16'h6463;
		end
		32'h0000FD92: begin
				q			<=			16'h6665;
		end
		32'h0000FD94: begin
				q			<=			16'h0000;
		end
		32'h0000FD96: begin
				q			<=			16'h0000;
		end
		32'h0000FD98: begin
				q			<=			16'h3130;
		end
		32'h0000FD9A: begin
				q			<=			16'h3332;
		end
		32'h0000FD9C: begin
				q			<=			16'h3534;
		end
		32'h0000FD9E: begin
				q			<=			16'h3736;
		end
		32'h0000FDA0: begin
				q			<=			16'h3938;
		end
		32'h0000FDA2: begin
				q			<=			16'h4241;
		end
		32'h0000FDA4: begin
				q			<=			16'h4443;
		end
		32'h0000FDA6: begin
				q			<=			16'h4645;
		end
		32'h0000FDA8: begin
				q			<=			16'h0000;
		end
		32'h0000FDAA: begin
				q			<=			16'h0000;
		end
		32'h0000FDAC: begin
				q			<=			16'h0030;
		end
		32'h0000FDAE: begin
				q			<=			16'h0000;
		end
		32'h0000FDB0: begin
				q			<=			16'h4E20;
		end
		32'h0000FDB2: begin
				q			<=			16'h4E61;
		end
		32'h0000FDB4: begin
				q			<=			16'h0020;
		end
		32'h0000FDB6: begin
				q			<=			16'h0000;
		end
		32'h0000FDB8: begin
				q			<=			16'h2D20;
		end
		32'h0000FDBA: begin
				q			<=			16'h6E49;
		end
		32'h0000FDBC: begin
				q			<=			16'h6966;
		end
		32'h0000FDBE: begin
				q			<=			16'h696E;
		end
		32'h0000FDC0: begin
				q			<=			16'h7974;
		end
		32'h0000FDC2: begin
				q			<=			16'h0020;
		end
		32'h0000FDC4: begin
				q			<=			16'h4920;
		end
		32'h0000FDC6: begin
				q			<=			16'h666E;
		end
		32'h0000FDC8: begin
				q			<=			16'h6E69;
		end
		32'h0000FDCA: begin
				q			<=			16'h7469;
		end
		32'h0000FDCC: begin
				q			<=			16'h2079;
		end
		32'h0000FDCE: begin
				q			<=			16'h0000;
		end
		32'h0000FDD0: begin
				q			<=			16'h614E;
		end
		32'h0000FDD2: begin
				q			<=			16'h004E;
		end
		32'h0000FDD4: begin
				q			<=			16'h2545;
		end
		32'h0000FDD6: begin
				q			<=			16'h0064;
		end
		32'h0000FDD8: begin
				q			<=			16'h0043;
		end
		32'h0000FDDA: begin
				q			<=			16'h0000;
		end
		32'h0000FDDC: begin
				q			<=			16'h4F50;
		end
		32'h0000FDDE: begin
				q			<=			16'h4953;
		end
		32'h0000FDE0: begin
				q			<=			16'h0058;
		end
		32'h0000FDE2: begin
				q			<=			16'h0000;
		end
		32'h0000FDE4: begin
				q			<=			16'h002E;
		end
		32'h0000FDE6: begin
				q			<=			16'h0000;
		end
		32'h0000FDE8: begin
				q			<=			16'h0010;
		end
		32'h0000FDEA: begin
				q			<=			16'h0000;
		end
		32'h0000FDEC: begin
				q			<=			16'h0000;
		end
		32'h0000FDEE: begin
				q			<=			16'h0000;
		end
		32'h0000FDF0: begin
				q			<=			16'h7A01;
		end
		32'h0000FDF2: begin
				q			<=			16'h0052;
		end
		32'h0000FDF4: begin
				q			<=			16'h7C01;
		end
		32'h0000FDF6: begin
				q			<=			16'h0105;
		end
		32'h0000FDF8: begin
				q			<=			16'h0D1B;
		end
		32'h0000FDFA: begin
				q			<=			16'h0002;
		end
		32'h0000FDFC: begin
				q			<=			16'h0048;
		end
		32'h0000FDFE: begin
				q			<=			16'h0000;
		end
		32'h0000FE00: begin
				q			<=			16'h0018;
		end
		32'h0000FE02: begin
				q			<=			16'h0000;
		end
		32'h0000FE04: begin
				q			<=			16'h2C38;
		end
		32'h0000FE06: begin
				q			<=			16'hFFFF;
		end
		32'h0000FE08: begin
				q			<=			16'h005C;
		end
		32'h0000FE0A: begin
				q			<=			16'h0000;
		end
		32'h0000FE0C: begin
				q			<=			16'h4400;
		end
		32'h0000FE0E: begin
				q			<=			16'h400E;
		end
		32'h0000FE10: begin
				q			<=			16'h9B48;
		end
		32'h0000FE12: begin
				q			<=			16'h440D;
		end
		32'h0000FE14: begin
				q			<=			16'h44DB;
		end
		32'h0000FE16: begin
				q			<=			16'h400E;
		end
		32'h0000FE18: begin
				q			<=			16'h9A48;
		end
		32'h0000FE1A: begin
				q			<=			16'h440C;
		end
		32'h0000FE1C: begin
				q			<=			16'h0B99;
		end
		32'h0000FE1E: begin
				q			<=			16'h9844;
		end
		32'h0000FE20: begin
				q			<=			16'h440A;
		end
		32'h0000FE22: begin
				q			<=			16'h0997;
		end
		32'h0000FE24: begin
				q			<=			16'hD744;
		end
		32'h0000FE26: begin
				q			<=			16'hD9D8;
		end
		32'h0000FE28: begin
				q			<=			16'hDBDA;
		end
		32'h0000FE2A: begin
				q			<=			16'h0E44;
		end
		32'h0000FE2C: begin
				q			<=			16'h4840;
		end
		32'h0000FE2E: begin
				q			<=			16'h0896;
		end
		32'h0000FE30: begin
				q			<=			16'h9544;
		end
		32'h0000FE32: begin
				q			<=			16'h4407;
		end
		32'h0000FE34: begin
				q			<=			16'h0694;
		end
		32'h0000FE36: begin
				q			<=			16'h9344;
		end
		32'h0000FE38: begin
				q			<=			16'h4405;
		end
		32'h0000FE3A: begin
				q			<=			16'h0492;
		end
		32'h0000FE3C: begin
				q			<=			16'h8944;
		end
		32'h0000FE3E: begin
				q			<=			16'h4403;
		end
		32'h0000FE40: begin
				q			<=			16'h0288;
		end
		32'h0000FE42: begin
				q			<=			16'h8144;
		end
		32'h0000FE44: begin
				q			<=			16'h0001;
		end
		32'h0000FE46: begin
				q			<=			16'h0000;
		end
		32'h0000FE48: begin
				q			<=			16'h001C;
		end
		32'h0000FE4A: begin
				q			<=			16'h0000;
		end
		32'h0000FE4C: begin
				q			<=			16'h0064;
		end
		32'h0000FE4E: begin
				q			<=			16'h0000;
		end
		32'h0000FE50: begin
				q			<=			16'h2C48;
		end
		32'h0000FE52: begin
				q			<=			16'hFFFF;
		end
		32'h0000FE54: begin
				q			<=			16'h0018;
		end
		32'h0000FE56: begin
				q			<=			16'h0000;
		end
		32'h0000FE58: begin
				q			<=			16'h4400;
		end
		32'h0000FE5A: begin
				q			<=			16'h100E;
		end
		32'h0000FE5C: begin
				q			<=			16'h8948;
		end
		32'h0000FE5E: begin
				q			<=			16'h4404;
		end
		32'h0000FE60: begin
				q			<=			16'h0288;
		end
		32'h0000FE62: begin
				q			<=			16'h8144;
		end
		32'h0000FE64: begin
				q			<=			16'h0001;
		end
		32'h0000FE66: begin
				q			<=			16'h0000;
		end
		32'h0000FE68: begin
				q			<=			16'h002C;
		end
		32'h0000FE6A: begin
				q			<=			16'h0000;
		end
		32'h0000FE6C: begin
				q			<=			16'h0000;
		end
		32'h0000FE6E: begin
				q			<=			16'h0000;
		end
		32'h0000FE70: begin
				q			<=			16'h7A01;
		end
		32'h0000FE72: begin
				q			<=			16'h0052;
		end
		32'h0000FE74: begin
				q			<=			16'h7C01;
		end
		32'h0000FE76: begin
				q			<=			16'h0101;
		end
		32'h0000FE78: begin
				q			<=			16'h0D1B;
		end
		32'h0000FE7A: begin
				q			<=			16'h0E02;
		end
		32'h0000FE7C: begin
				q			<=			16'h9B40;
		end
		32'h0000FE7E: begin
				q			<=			16'h9A0D;
		end
		32'h0000FE80: begin
				q			<=			16'h990C;
		end
		32'h0000FE82: begin
				q			<=			16'h980B;
		end
		32'h0000FE84: begin
				q			<=			16'h970A;
		end
		32'h0000FE86: begin
				q			<=			16'h9609;
		end
		32'h0000FE88: begin
				q			<=			16'h9508;
		end
		32'h0000FE8A: begin
				q			<=			16'h9407;
		end
		32'h0000FE8C: begin
				q			<=			16'h9306;
		end
		32'h0000FE8E: begin
				q			<=			16'h9205;
		end
		32'h0000FE90: begin
				q			<=			16'h8904;
		end
		32'h0000FE92: begin
				q			<=			16'h8803;
		end
		32'h0000FE94: begin
				q			<=			16'h8102;
		end
		32'h0000FE96: begin
				q			<=			16'h0001;
		end
		32'h0000FE98: begin
				q			<=			16'h0044;
		end
		32'h0000FE9A: begin
				q			<=			16'h0000;
		end
		32'h0000FE9C: begin
				q			<=			16'h0034;
		end
		32'h0000FE9E: begin
				q			<=			16'h0000;
		end
		32'h0000FEA0: begin
				q			<=			16'h2C10;
		end
		32'h0000FEA2: begin
				q			<=			16'hFFFF;
		end
		32'h0000FEA4: begin
				q			<=			16'h0048;
		end
		32'h0000FEA6: begin
				q			<=			16'h0000;
		end
		32'h0000FEA8: begin
				q			<=			16'h4400;
		end
		32'h0000FEAA: begin
				q			<=			16'h44DB;
		end
		32'h0000FEAC: begin
				q			<=			16'h0EDB;
		end
		32'h0000FEAE: begin
				q			<=			16'h4430;
		end
		32'h0000FEB0: begin
				q			<=			16'h44DA;
		end
		32'h0000FEB2: begin
				q			<=			16'h44D9;
		end
		32'h0000FEB4: begin
				q			<=			16'h44D8;
		end
		32'h0000FEB6: begin
				q			<=			16'h44D7;
		end
		32'h0000FEB8: begin
				q			<=			16'hD8D7;
		end
		32'h0000FEBA: begin
				q			<=			16'hDAD9;
		end
		32'h0000FEBC: begin
				q			<=			16'h0EDB;
		end
		32'h0000FEBE: begin
				q			<=			16'h4420;
		end
		32'h0000FEC0: begin
				q			<=			16'h44D6;
		end
		32'h0000FEC2: begin
				q			<=			16'h44D5;
		end
		32'h0000FEC4: begin
				q			<=			16'h44D4;
		end
		32'h0000FEC6: begin
				q			<=			16'h44D3;
		end
		32'h0000FEC8: begin
				q			<=			16'hD4D3;
		end
		32'h0000FECA: begin
				q			<=			16'hD6D5;
		end
		32'h0000FECC: begin
				q			<=			16'hD9D8;
		end
		32'h0000FECE: begin
				q			<=			16'hDBDA;
		end
		32'h0000FED0: begin
				q			<=			16'h100E;
		end
		32'h0000FED2: begin
				q			<=			16'hD244;
		end
		32'h0000FED4: begin
				q			<=			16'hC944;
		end
		32'h0000FED6: begin
				q			<=			16'hC844;
		end
		32'h0000FED8: begin
				q			<=			16'hC144;
		end
		32'h0000FEDA: begin
				q			<=			16'h0E44;
		end
		32'h0000FEDC: begin
				q			<=			16'h0000;
		end
		32'h0000FEDE: begin
				q			<=			16'h0000;
		end
		32'h0000FEE0: begin
				q			<=			16'h0010;
		end
		32'h0000FEE2: begin
				q			<=			16'h0000;
		end
		32'h0000FEE4: begin
				q			<=			16'h0000;
		end
		32'h0000FEE6: begin
				q			<=			16'h0000;
		end
		32'h0000FEE8: begin
				q			<=			16'h7A01;
		end
		32'h0000FEEA: begin
				q			<=			16'h0052;
		end
		32'h0000FEEC: begin
				q			<=			16'h7C01;
		end
		32'h0000FEEE: begin
				q			<=			16'h0101;
		end
		32'h0000FEF0: begin
				q			<=			16'h0D1B;
		end
		32'h0000FEF2: begin
				q			<=			16'h0002;
		end
		32'h0000FEF4: begin
				q			<=			16'h0010;
		end
		32'h0000FEF6: begin
				q			<=			16'h0000;
		end
		32'h0000FEF8: begin
				q			<=			16'h0018;
		end
		32'h0000FEFA: begin
				q			<=			16'h0000;
		end
		32'h0000FEFC: begin
				q			<=			16'hABB0;
		end
		32'h0000FEFE: begin
				q			<=			16'hFFFF;
		end
		32'h0000FF00: begin
				q			<=			16'h0434;
		end
		32'h0000FF02: begin
				q			<=			16'h0000;
		end
		32'h0000FF04: begin
				q			<=			16'h0000;
		end
		32'h0000FF06: begin
				q			<=			16'h0000;
		end
		32'h0000FF08: begin
				q			<=			16'h0010;
		end
		32'h0000FF0A: begin
				q			<=			16'h0000;
		end
		32'h0000FF0C: begin
				q			<=			16'h002C;
		end
		32'h0000FF0E: begin
				q			<=			16'h0000;
		end
		32'h0000FF10: begin
				q			<=			16'hAFD4;
		end
		32'h0000FF12: begin
				q			<=			16'hFFFF;
		end
		32'h0000FF14: begin
				q			<=			16'h0410;
		end
		32'h0000FF16: begin
				q			<=			16'h0000;
		end
		32'h0000FF18: begin
				q			<=			16'h0000;
		end
		32'h0000FF1A: begin
				q			<=			16'h0000;
		end
		32'h0000FF1C: begin
				q			<=			16'h0000;
		end
		32'h0000FF1E: begin
				q			<=			16'h0000;
		end
		32'h0000FF20: begin
				q			<=			16'h0000;
		end
		32'h0000FF22: begin
				q			<=			16'h0000;
		end
		32'h0000FF24: begin
				q			<=			16'h0000;
		end
		32'h0000FF26: begin
				q			<=			16'h3FF0;
		end
		32'h0000FF28: begin
				q			<=			16'h0000;
		end
		32'h0000FF2A: begin
				q			<=			16'h0000;
		end
		32'h0000FF2C: begin
				q			<=			16'h0000;
		end
		32'h0000FF2E: begin
				q			<=			16'h4024;
		end
		32'h0000FF30: begin
				q			<=			16'h0000;
		end
		32'h0000FF32: begin
				q			<=			16'h0000;
		end
		32'h0000FF34: begin
				q			<=			16'h0000;
		end
		32'h0000FF36: begin
				q			<=			16'h4350;
		end
		32'h0000FF38: begin
				q			<=			16'h0000;
		end
		32'h0000FF3A: begin
				q			<=			16'h0000;
		end
		32'h0000FF3C: begin
				q			<=			16'h0224;
		end
		32'h0000FF3E: begin
				q			<=			16'h0001;
		end
		32'h0000FF40: begin
				q			<=			16'h028C;
		end
		32'h0000FF42: begin
				q			<=			16'h0001;
		end
		32'h0000FF44: begin
				q			<=			16'h02F4;
		end
		32'h0000FF46: begin
				q			<=			16'h0001;
		end
		32'h0000FF48: begin
				q			<=			16'h0000;
		end
		32'h0000FF4A: begin
				q			<=			16'h0000;
		end
		32'h0000FF4C: begin
				q			<=			16'h0000;
		end
		32'h0000FF4E: begin
				q			<=			16'h0000;
		end
		32'h0000FF50: begin
				q			<=			16'h0000;
		end
		32'h0000FF52: begin
				q			<=			16'h0000;
		end
		32'h0000FF54: begin
				q			<=			16'h0000;
		end
		32'h0000FF56: begin
				q			<=			16'h0000;
		end
		32'h0000FF58: begin
				q			<=			16'h0000;
		end
		32'h0000FF5A: begin
				q			<=			16'h0000;
		end
		32'h0000FF5C: begin
				q			<=			16'h0000;
		end
		32'h0000FF5E: begin
				q			<=			16'h0000;
		end
		32'h0000FF60: begin
				q			<=			16'h0000;
		end
		32'h0000FF62: begin
				q			<=			16'h0000;
		end
		32'h0000FF64: begin
				q			<=			16'h0000;
		end
		32'h0000FF66: begin
				q			<=			16'h0000;
		end
		32'h0000FF68: begin
				q			<=			16'h0000;
		end
		32'h0000FF6A: begin
				q			<=			16'h0000;
		end
		32'h0000FF6C: begin
				q			<=			16'h0000;
		end
		32'h0000FF6E: begin
				q			<=			16'h0000;
		end
		32'h0000FF70: begin
				q			<=			16'h0000;
		end
		32'h0000FF72: begin
				q			<=			16'h0000;
		end
		32'h0000FF74: begin
				q			<=			16'h0000;
		end
		32'h0000FF76: begin
				q			<=			16'h0000;
		end
		32'h0000FF78: begin
				q			<=			16'h0000;
		end
		32'h0000FF7A: begin
				q			<=			16'h0000;
		end
		32'h0000FF7C: begin
				q			<=			16'h0000;
		end
		32'h0000FF7E: begin
				q			<=			16'h0000;
		end
		32'h0000FF80: begin
				q			<=			16'h0000;
		end
		32'h0000FF82: begin
				q			<=			16'h0000;
		end
		32'h0000FF84: begin
				q			<=			16'h0000;
		end
		32'h0000FF86: begin
				q			<=			16'h0000;
		end
		32'h0000FF88: begin
				q			<=			16'h0000;
		end
		32'h0000FF8A: begin
				q			<=			16'h0000;
		end
		32'h0000FF8C: begin
				q			<=			16'h0000;
		end
		32'h0000FF8E: begin
				q			<=			16'h0000;
		end
		32'h0000FF90: begin
				q			<=			16'h0000;
		end
		32'h0000FF92: begin
				q			<=			16'h0000;
		end
		32'h0000FF94: begin
				q			<=			16'h0000;
		end
		32'h0000FF96: begin
				q			<=			16'h0000;
		end
		32'h0000FF98: begin
				q			<=			16'h0000;
		end
		32'h0000FF9A: begin
				q			<=			16'h0000;
		end
		32'h0000FF9C: begin
				q			<=			16'h0000;
		end
		32'h0000FF9E: begin
				q			<=			16'h0000;
		end
		32'h0000FFA0: begin
				q			<=			16'h0000;
		end
		32'h0000FFA2: begin
				q			<=			16'h0000;
		end
		32'h0000FFA4: begin
				q			<=			16'h0000;
		end
		32'h0000FFA6: begin
				q			<=			16'h0000;
		end
		32'h0000FFA8: begin
				q			<=			16'h0000;
		end
		32'h0000FFAA: begin
				q			<=			16'h0000;
		end
		32'h0000FFAC: begin
				q			<=			16'h0000;
		end
		32'h0000FFAE: begin
				q			<=			16'h0000;
		end
		32'h0000FFB0: begin
				q			<=			16'h0000;
		end
		32'h0000FFB2: begin
				q			<=			16'h0000;
		end
		32'h0000FFB4: begin
				q			<=			16'h0000;
		end
		32'h0000FFB6: begin
				q			<=			16'h0000;
		end
		32'h0000FFB8: begin
				q			<=			16'h0000;
		end
		32'h0000FFBA: begin
				q			<=			16'h0000;
		end
		32'h0000FFBC: begin
				q			<=			16'h0000;
		end
		32'h0000FFBE: begin
				q			<=			16'h0000;
		end
		32'h0000FFC0: begin
				q			<=			16'h0000;
		end
		32'h0000FFC2: begin
				q			<=			16'h0000;
		end
		32'h0000FFC4: begin
				q			<=			16'h0000;
		end
		32'h0000FFC6: begin
				q			<=			16'h0000;
		end
		32'h0000FFC8: begin
				q			<=			16'h0000;
		end
		32'h0000FFCA: begin
				q			<=			16'h0000;
		end
		32'h0000FFCC: begin
				q			<=			16'h0000;
		end
		32'h0000FFCE: begin
				q			<=			16'h0000;
		end
		32'h0000FFD0: begin
				q			<=			16'h0000;
		end
		32'h0000FFD2: begin
				q			<=			16'h0000;
		end
		32'h0000FFD4: begin
				q			<=			16'h0000;
		end
		32'h0000FFD6: begin
				q			<=			16'h0000;
		end
		32'h0000FFD8: begin
				q			<=			16'h0000;
		end
		32'h0000FFDA: begin
				q			<=			16'h0000;
		end
		32'h0000FFDC: begin
				q			<=			16'h0000;
		end
		32'h0000FFDE: begin
				q			<=			16'h0000;
		end
		32'h0000FFE0: begin
				q			<=			16'h0001;
		end
		32'h0000FFE2: begin
				q			<=			16'h0000;
		end
		32'h0000FFE4: begin
				q			<=			16'h0000;
		end
		32'h0000FFE6: begin
				q			<=			16'h0000;
		end
		32'h0000FFE8: begin
				q			<=			16'h330E;
		end
		32'h0000FFEA: begin
				q			<=			16'hABCD;
		end
		32'h0000FFEC: begin
				q			<=			16'h1234;
		end
		32'h0000FFEE: begin
				q			<=			16'hE66D;
		end
		32'h0000FFF0: begin
				q			<=			16'hDEEC;
		end
		32'h0000FFF2: begin
				q			<=			16'h0005;
		end
		32'h0000FFF4: begin
				q			<=			16'h000B;
		end
		32'h0000FFF6: begin
				q			<=			16'h0000;
		end
		32'h0000FFF8: begin
				q			<=			16'h0000;
		end
		32'h0000FFFA: begin
				q			<=			16'h0000;
		end
		32'h0000FFFC: begin
				q			<=			16'h0000;
		end
		32'h0000FFFE: begin
				q			<=			16'h0000;
		end
		32'h00010000: begin
				q			<=			16'h0000;
		end
		32'h00010002: begin
				q			<=			16'h0000;
		end
		32'h00010004: begin
				q			<=			16'h0000;
		end
		32'h00010006: begin
				q			<=			16'h0000;
		end
		32'h00010008: begin
				q			<=			16'h0000;
		end
		32'h0001000A: begin
				q			<=			16'h0000;
		end
		32'h0001000C: begin
				q			<=			16'h0000;
		end
		32'h0001000E: begin
				q			<=			16'h0000;
		end
		32'h00010010: begin
				q			<=			16'h0000;
		end
		32'h00010012: begin
				q			<=			16'h0000;
		end
		32'h00010014: begin
				q			<=			16'h0000;
		end
		32'h00010016: begin
				q			<=			16'h0000;
		end
		32'h00010018: begin
				q			<=			16'h0000;
		end
		32'h0001001A: begin
				q			<=			16'h0000;
		end
		32'h0001001C: begin
				q			<=			16'h0000;
		end
		32'h0001001E: begin
				q			<=			16'h0000;
		end
		32'h00010020: begin
				q			<=			16'h0000;
		end
		32'h00010022: begin
				q			<=			16'h0000;
		end
		32'h00010024: begin
				q			<=			16'h0000;
		end
		32'h00010026: begin
				q			<=			16'h0000;
		end
		32'h00010028: begin
				q			<=			16'h0000;
		end
		32'h0001002A: begin
				q			<=			16'h0000;
		end
		32'h0001002C: begin
				q			<=			16'h0000;
		end
		32'h0001002E: begin
				q			<=			16'h0000;
		end
		32'h00010030: begin
				q			<=			16'h0000;
		end
		32'h00010032: begin
				q			<=			16'h0000;
		end
		32'h00010034: begin
				q			<=			16'h0000;
		end
		32'h00010036: begin
				q			<=			16'h0000;
		end
		32'h00010038: begin
				q			<=			16'h0000;
		end
		32'h0001003A: begin
				q			<=			16'h0000;
		end
		32'h0001003C: begin
				q			<=			16'h0000;
		end
		32'h0001003E: begin
				q			<=			16'h0000;
		end
		32'h00010040: begin
				q			<=			16'h0000;
		end
		32'h00010042: begin
				q			<=			16'h0000;
		end
		32'h00010044: begin
				q			<=			16'h0000;
		end
		32'h00010046: begin
				q			<=			16'h0000;
		end
		32'h00010048: begin
				q			<=			16'h0000;
		end
		32'h0001004A: begin
				q			<=			16'h0000;
		end
		32'h0001004C: begin
				q			<=			16'h0000;
		end
		32'h0001004E: begin
				q			<=			16'h0000;
		end
		32'h00010050: begin
				q			<=			16'h0000;
		end
		32'h00010052: begin
				q			<=			16'h0000;
		end
		32'h00010054: begin
				q			<=			16'h0000;
		end
		32'h00010056: begin
				q			<=			16'h0000;
		end
		32'h00010058: begin
				q			<=			16'h0000;
		end
		32'h0001005A: begin
				q			<=			16'h0000;
		end
		32'h0001005C: begin
				q			<=			16'h0000;
		end
		32'h0001005E: begin
				q			<=			16'h0000;
		end
		32'h00010060: begin
				q			<=			16'h0000;
		end
		32'h00010062: begin
				q			<=			16'h0000;
		end
		32'h00010064: begin
				q			<=			16'h0000;
		end
		32'h00010066: begin
				q			<=			16'h0000;
		end
		32'h00010068: begin
				q			<=			16'h0000;
		end
		32'h0001006A: begin
				q			<=			16'h0000;
		end
		32'h0001006C: begin
				q			<=			16'h0000;
		end
		32'h0001006E: begin
				q			<=			16'h0000;
		end
		32'h00010070: begin
				q			<=			16'h0000;
		end
		32'h00010072: begin
				q			<=			16'h0000;
		end
		32'h00010074: begin
				q			<=			16'h0000;
		end
		32'h00010076: begin
				q			<=			16'h0000;
		end
		32'h00010078: begin
				q			<=			16'h0000;
		end
		32'h0001007A: begin
				q			<=			16'h0000;
		end
		32'h0001007C: begin
				q			<=			16'h0000;
		end
		32'h0001007E: begin
				q			<=			16'h0000;
		end
		32'h00010080: begin
				q			<=			16'h0000;
		end
		32'h00010082: begin
				q			<=			16'h0000;
		end
		32'h00010084: begin
				q			<=			16'h0000;
		end
		32'h00010086: begin
				q			<=			16'h0000;
		end
		32'h00010088: begin
				q			<=			16'h0000;
		end
		32'h0001008A: begin
				q			<=			16'h0000;
		end
		32'h0001008C: begin
				q			<=			16'h0000;
		end
		32'h0001008E: begin
				q			<=			16'h0000;
		end
		32'h00010090: begin
				q			<=			16'h0000;
		end
		32'h00010092: begin
				q			<=			16'h0000;
		end
		32'h00010094: begin
				q			<=			16'h0000;
		end
		32'h00010096: begin
				q			<=			16'h0000;
		end
		32'h00010098: begin
				q			<=			16'h0000;
		end
		32'h0001009A: begin
				q			<=			16'h0000;
		end
		32'h0001009C: begin
				q			<=			16'h0000;
		end
		32'h0001009E: begin
				q			<=			16'h0000;
		end
		32'h000100A0: begin
				q			<=			16'h0000;
		end
		32'h000100A2: begin
				q			<=			16'h0000;
		end
		32'h000100A4: begin
				q			<=			16'h0000;
		end
		32'h000100A6: begin
				q			<=			16'h0000;
		end
		32'h000100A8: begin
				q			<=			16'h0000;
		end
		32'h000100AA: begin
				q			<=			16'h0000;
		end
		32'h000100AC: begin
				q			<=			16'h0000;
		end
		32'h000100AE: begin
				q			<=			16'h0000;
		end
		32'h000100B0: begin
				q			<=			16'h0000;
		end
		32'h000100B2: begin
				q			<=			16'h0000;
		end
		32'h000100B4: begin
				q			<=			16'h0000;
		end
		32'h000100B6: begin
				q			<=			16'h0000;
		end
		32'h000100B8: begin
				q			<=			16'h0000;
		end
		32'h000100BA: begin
				q			<=			16'h0000;
		end
		32'h000100BC: begin
				q			<=			16'h0000;
		end
		32'h000100BE: begin
				q			<=			16'h0000;
		end
		32'h000100C0: begin
				q			<=			16'h0000;
		end
		32'h000100C2: begin
				q			<=			16'h0000;
		end
		32'h000100C4: begin
				q			<=			16'h0000;
		end
		32'h000100C6: begin
				q			<=			16'h0000;
		end
		32'h000100C8: begin
				q			<=			16'h0000;
		end
		32'h000100CA: begin
				q			<=			16'h0000;
		end
		32'h000100CC: begin
				q			<=			16'h0000;
		end
		32'h000100CE: begin
				q			<=			16'h0000;
		end
		32'h000100D0: begin
				q			<=			16'h0000;
		end
		32'h000100D2: begin
				q			<=			16'h0000;
		end
		32'h000100D4: begin
				q			<=			16'h0000;
		end
		32'h000100D6: begin
				q			<=			16'h0000;
		end
		32'h000100D8: begin
				q			<=			16'h0000;
		end
		32'h000100DA: begin
				q			<=			16'h0000;
		end
		32'h000100DC: begin
				q			<=			16'h0000;
		end
		32'h000100DE: begin
				q			<=			16'h0000;
		end
		32'h000100E0: begin
				q			<=			16'h0000;
		end
		32'h000100E2: begin
				q			<=			16'h0000;
		end
		32'h000100E4: begin
				q			<=			16'h0000;
		end
		32'h000100E6: begin
				q			<=			16'h0000;
		end
		32'h000100E8: begin
				q			<=			16'h0000;
		end
		32'h000100EA: begin
				q			<=			16'h0000;
		end
		32'h000100EC: begin
				q			<=			16'h0000;
		end
		32'h000100EE: begin
				q			<=			16'h0000;
		end
		32'h000100F0: begin
				q			<=			16'h0000;
		end
		32'h000100F2: begin
				q			<=			16'h0000;
		end
		32'h000100F4: begin
				q			<=			16'h0000;
		end
		32'h000100F6: begin
				q			<=			16'h0000;
		end
		32'h000100F8: begin
				q			<=			16'h0000;
		end
		32'h000100FA: begin
				q			<=			16'h0000;
		end
		32'h000100FC: begin
				q			<=			16'h0000;
		end
		32'h000100FE: begin
				q			<=			16'h0000;
		end
		32'h00010100: begin
				q			<=			16'h0000;
		end
		32'h00010102: begin
				q			<=			16'h0000;
		end
		32'h00010104: begin
				q			<=			16'h0000;
		end
		32'h00010106: begin
				q			<=			16'h0000;
		end
		32'h00010108: begin
				q			<=			16'h0000;
		end
		32'h0001010A: begin
				q			<=			16'h0000;
		end
		32'h0001010C: begin
				q			<=			16'h0000;
		end
		32'h0001010E: begin
				q			<=			16'h0000;
		end
		32'h00010110: begin
				q			<=			16'h0000;
		end
		32'h00010112: begin
				q			<=			16'h0000;
		end
		32'h00010114: begin
				q			<=			16'h0000;
		end
		32'h00010116: begin
				q			<=			16'h0000;
		end
		32'h00010118: begin
				q			<=			16'h0000;
		end
		32'h0001011A: begin
				q			<=			16'h0000;
		end
		32'h0001011C: begin
				q			<=			16'h0000;
		end
		32'h0001011E: begin
				q			<=			16'h0000;
		end
		32'h00010120: begin
				q			<=			16'h0000;
		end
		32'h00010122: begin
				q			<=			16'h0000;
		end
		32'h00010124: begin
				q			<=			16'h0000;
		end
		32'h00010126: begin
				q			<=			16'h0000;
		end
		32'h00010128: begin
				q			<=			16'h0000;
		end
		32'h0001012A: begin
				q			<=			16'h0000;
		end
		32'h0001012C: begin
				q			<=			16'h0000;
		end
		32'h0001012E: begin
				q			<=			16'h0000;
		end
		32'h00010130: begin
				q			<=			16'h0000;
		end
		32'h00010132: begin
				q			<=			16'h0000;
		end
		32'h00010134: begin
				q			<=			16'h0000;
		end
		32'h00010136: begin
				q			<=			16'h0000;
		end
		32'h00010138: begin
				q			<=			16'h0000;
		end
		32'h0001013A: begin
				q			<=			16'h0000;
		end
		32'h0001013C: begin
				q			<=			16'h0000;
		end
		32'h0001013E: begin
				q			<=			16'h0000;
		end
		32'h00010140: begin
				q			<=			16'h0000;
		end
		32'h00010142: begin
				q			<=			16'h0000;
		end
		32'h00010144: begin
				q			<=			16'h0000;
		end
		32'h00010146: begin
				q			<=			16'h0000;
		end
		32'h00010148: begin
				q			<=			16'h0000;
		end
		32'h0001014A: begin
				q			<=			16'h0000;
		end
		32'h0001014C: begin
				q			<=			16'h0000;
		end
		32'h0001014E: begin
				q			<=			16'h0000;
		end
		32'h00010150: begin
				q			<=			16'h0000;
		end
		32'h00010152: begin
				q			<=			16'h0000;
		end
		32'h00010154: begin
				q			<=			16'h0000;
		end
		32'h00010156: begin
				q			<=			16'h0000;
		end
		32'h00010158: begin
				q			<=			16'h0000;
		end
		32'h0001015A: begin
				q			<=			16'h0000;
		end
		32'h0001015C: begin
				q			<=			16'h0000;
		end
		32'h0001015E: begin
				q			<=			16'h0000;
		end
		32'h00010160: begin
				q			<=			16'h0000;
		end
		32'h00010162: begin
				q			<=			16'h0000;
		end
		32'h00010164: begin
				q			<=			16'h0000;
		end
		32'h00010166: begin
				q			<=			16'h0000;
		end
		32'h00010168: begin
				q			<=			16'h0000;
		end
		32'h0001016A: begin
				q			<=			16'h0000;
		end
		32'h0001016C: begin
				q			<=			16'h0000;
		end
		32'h0001016E: begin
				q			<=			16'h0000;
		end
		32'h00010170: begin
				q			<=			16'h0000;
		end
		32'h00010172: begin
				q			<=			16'h0000;
		end
		32'h00010174: begin
				q			<=			16'h0000;
		end
		32'h00010176: begin
				q			<=			16'h0000;
		end
		32'h00010178: begin
				q			<=			16'h0000;
		end
		32'h0001017A: begin
				q			<=			16'h0000;
		end
		32'h0001017C: begin
				q			<=			16'h0000;
		end
		32'h0001017E: begin
				q			<=			16'h0000;
		end
		32'h00010180: begin
				q			<=			16'h0000;
		end
		32'h00010182: begin
				q			<=			16'h0000;
		end
		32'h00010184: begin
				q			<=			16'h0000;
		end
		32'h00010186: begin
				q			<=			16'h0000;
		end
		32'h00010188: begin
				q			<=			16'h0000;
		end
		32'h0001018A: begin
				q			<=			16'h0000;
		end
		32'h0001018C: begin
				q			<=			16'h0000;
		end
		32'h0001018E: begin
				q			<=			16'h0000;
		end
		32'h00010190: begin
				q			<=			16'h0000;
		end
		32'h00010192: begin
				q			<=			16'h0000;
		end
		32'h00010194: begin
				q			<=			16'h0000;
		end
		32'h00010196: begin
				q			<=			16'h0000;
		end
		32'h00010198: begin
				q			<=			16'h0000;
		end
		32'h0001019A: begin
				q			<=			16'h0000;
		end
		32'h0001019C: begin
				q			<=			16'h0000;
		end
		32'h0001019E: begin
				q			<=			16'h0000;
		end
		32'h000101A0: begin
				q			<=			16'h0000;
		end
		32'h000101A2: begin
				q			<=			16'h0000;
		end
		32'h000101A4: begin
				q			<=			16'h0000;
		end
		32'h000101A6: begin
				q			<=			16'h0000;
		end
		32'h000101A8: begin
				q			<=			16'h0000;
		end
		32'h000101AA: begin
				q			<=			16'h0000;
		end
		32'h000101AC: begin
				q			<=			16'h0000;
		end
		32'h000101AE: begin
				q			<=			16'h0000;
		end
		32'h000101B0: begin
				q			<=			16'h0000;
		end
		32'h000101B2: begin
				q			<=			16'h0000;
		end
		32'h000101B4: begin
				q			<=			16'h0000;
		end
		32'h000101B6: begin
				q			<=			16'h0000;
		end
		32'h000101B8: begin
				q			<=			16'h0000;
		end
		32'h000101BA: begin
				q			<=			16'h0000;
		end
		32'h000101BC: begin
				q			<=			16'h0000;
		end
		32'h000101BE: begin
				q			<=			16'h0000;
		end
		32'h000101C0: begin
				q			<=			16'h0000;
		end
		32'h000101C2: begin
				q			<=			16'h0000;
		end
		32'h000101C4: begin
				q			<=			16'h0000;
		end
		32'h000101C6: begin
				q			<=			16'h0000;
		end
		32'h000101C8: begin
				q			<=			16'h0000;
		end
		32'h000101CA: begin
				q			<=			16'h0000;
		end
		32'h000101CC: begin
				q			<=			16'h0000;
		end
		32'h000101CE: begin
				q			<=			16'h0000;
		end
		32'h000101D0: begin
				q			<=			16'h0000;
		end
		32'h000101D2: begin
				q			<=			16'h0000;
		end
		32'h000101D4: begin
				q			<=			16'h0000;
		end
		32'h000101D6: begin
				q			<=			16'h0000;
		end
		32'h000101D8: begin
				q			<=			16'h0000;
		end
		32'h000101DA: begin
				q			<=			16'h0000;
		end
		32'h000101DC: begin
				q			<=			16'h0000;
		end
		32'h000101DE: begin
				q			<=			16'h0000;
		end
		32'h000101E0: begin
				q			<=			16'h0000;
		end
		32'h000101E2: begin
				q			<=			16'h0000;
		end
		32'h000101E4: begin
				q			<=			16'h0000;
		end
		32'h000101E6: begin
				q			<=			16'h0000;
		end
		32'h000101E8: begin
				q			<=			16'h0000;
		end
		32'h000101EA: begin
				q			<=			16'h0000;
		end
		32'h000101EC: begin
				q			<=			16'h0000;
		end
		32'h000101EE: begin
				q			<=			16'h0000;
		end
		32'h000101F0: begin
				q			<=			16'h0000;
		end
		32'h000101F2: begin
				q			<=			16'h0000;
		end
		32'h000101F4: begin
				q			<=			16'h0000;
		end
		32'h000101F6: begin
				q			<=			16'h0000;
		end
		32'h000101F8: begin
				q			<=			16'h0000;
		end
		32'h000101FA: begin
				q			<=			16'h0000;
		end
		32'h000101FC: begin
				q			<=			16'h0000;
		end
		32'h000101FE: begin
				q			<=			16'h0000;
		end
		32'h00010200: begin
				q			<=			16'h0000;
		end
		32'h00010202: begin
				q			<=			16'h0000;
		end
		32'h00010204: begin
				q			<=			16'h0000;
		end
		32'h00010206: begin
				q			<=			16'h0000;
		end
		32'h00010208: begin
				q			<=			16'h0000;
		end
		32'h0001020A: begin
				q			<=			16'h0000;
		end
		32'h0001020C: begin
				q			<=			16'h0000;
		end
		32'h0001020E: begin
				q			<=			16'h0000;
		end
		32'h00010210: begin
				q			<=			16'h0000;
		end
		32'h00010212: begin
				q			<=			16'h0000;
		end
		32'h00010214: begin
				q			<=			16'h0000;
		end
		32'h00010216: begin
				q			<=			16'h0000;
		end
		32'h00010218: begin
				q			<=			16'h0000;
		end
		32'h0001021A: begin
				q			<=			16'h0000;
		end
		32'h0001021C: begin
				q			<=			16'h0000;
		end
		32'h0001021E: begin
				q			<=			16'h0000;
		end
		32'h00010220: begin
				q			<=			16'h0000;
		end
		32'h00010222: begin
				q			<=			16'h0000;
		end
		32'h00010224: begin
				q			<=			16'h0000;
		end
		32'h00010226: begin
				q			<=			16'h0000;
		end
		32'h00010228: begin
				q			<=			16'h0000;
		end
		32'h0001022A: begin
				q			<=			16'h0000;
		end
		32'h0001022C: begin
				q			<=			16'h0000;
		end
		32'h0001022E: begin
				q			<=			16'h0000;
		end
		32'h00010230: begin
				q			<=			16'h0000;
		end
		32'h00010232: begin
				q			<=			16'h0000;
		end
		32'h00010234: begin
				q			<=			16'h0000;
		end
		32'h00010236: begin
				q			<=			16'h0000;
		end
		32'h00010238: begin
				q			<=			16'h0000;
		end
		32'h0001023A: begin
				q			<=			16'h0000;
		end
		32'h0001023C: begin
				q			<=			16'h0000;
		end
		32'h0001023E: begin
				q			<=			16'h0000;
		end
		32'h00010240: begin
				q			<=			16'h0000;
		end
		32'h00010242: begin
				q			<=			16'h0000;
		end
		32'h00010244: begin
				q			<=			16'h0000;
		end
		32'h00010246: begin
				q			<=			16'h0000;
		end
		32'h00010248: begin
				q			<=			16'h0000;
		end
		32'h0001024A: begin
				q			<=			16'h0000;
		end
		32'h0001024C: begin
				q			<=			16'h0000;
		end
		32'h0001024E: begin
				q			<=			16'h0000;
		end
		32'h00010250: begin
				q			<=			16'h0000;
		end
		32'h00010252: begin
				q			<=			16'h0000;
		end
		32'h00010254: begin
				q			<=			16'h0000;
		end
		32'h00010256: begin
				q			<=			16'h0000;
		end
		32'h00010258: begin
				q			<=			16'h0000;
		end
		32'h0001025A: begin
				q			<=			16'h0000;
		end
		32'h0001025C: begin
				q			<=			16'h0000;
		end
		32'h0001025E: begin
				q			<=			16'h0000;
		end
		32'h00010260: begin
				q			<=			16'h0000;
		end
		32'h00010262: begin
				q			<=			16'h0000;
		end
		32'h00010264: begin
				q			<=			16'h0000;
		end
		32'h00010266: begin
				q			<=			16'h0000;
		end
		32'h00010268: begin
				q			<=			16'h0000;
		end
		32'h0001026A: begin
				q			<=			16'h0000;
		end
		32'h0001026C: begin
				q			<=			16'h0000;
		end
		32'h0001026E: begin
				q			<=			16'h0000;
		end
		32'h00010270: begin
				q			<=			16'h0000;
		end
		32'h00010272: begin
				q			<=			16'h0000;
		end
		32'h00010274: begin
				q			<=			16'h0000;
		end
		32'h00010276: begin
				q			<=			16'h0000;
		end
		32'h00010278: begin
				q			<=			16'h0000;
		end
		32'h0001027A: begin
				q			<=			16'h0000;
		end
		32'h0001027C: begin
				q			<=			16'h0000;
		end
		32'h0001027E: begin
				q			<=			16'h0000;
		end
		32'h00010280: begin
				q			<=			16'h0000;
		end
		32'h00010282: begin
				q			<=			16'h0000;
		end
		32'h00010284: begin
				q			<=			16'h0000;
		end
		32'h00010286: begin
				q			<=			16'h0000;
		end
		32'h00010288: begin
				q			<=			16'h0000;
		end
		32'h0001028A: begin
				q			<=			16'h0000;
		end
		32'h0001028C: begin
				q			<=			16'h0000;
		end
		32'h0001028E: begin
				q			<=			16'h0000;
		end
		32'h00010290: begin
				q			<=			16'h0000;
		end
		32'h00010292: begin
				q			<=			16'h0000;
		end
		32'h00010294: begin
				q			<=			16'h0000;
		end
		32'h00010296: begin
				q			<=			16'h0000;
		end
		32'h00010298: begin
				q			<=			16'h0000;
		end
		32'h0001029A: begin
				q			<=			16'h0000;
		end
		32'h0001029C: begin
				q			<=			16'h0000;
		end
		32'h0001029E: begin
				q			<=			16'h0000;
		end
		32'h000102A0: begin
				q			<=			16'h0000;
		end
		32'h000102A2: begin
				q			<=			16'h0000;
		end
		32'h000102A4: begin
				q			<=			16'h0000;
		end
		32'h000102A6: begin
				q			<=			16'h0000;
		end
		32'h000102A8: begin
				q			<=			16'h0000;
		end
		32'h000102AA: begin
				q			<=			16'h0000;
		end
		32'h000102AC: begin
				q			<=			16'h0000;
		end
		32'h000102AE: begin
				q			<=			16'h0000;
		end
		32'h000102B0: begin
				q			<=			16'h0000;
		end
		32'h000102B2: begin
				q			<=			16'h0000;
		end
		32'h000102B4: begin
				q			<=			16'h0000;
		end
		32'h000102B6: begin
				q			<=			16'h0000;
		end
		32'h000102B8: begin
				q			<=			16'h0000;
		end
		32'h000102BA: begin
				q			<=			16'h0000;
		end
		32'h000102BC: begin
				q			<=			16'h0000;
		end
		32'h000102BE: begin
				q			<=			16'h0000;
		end
		32'h000102C0: begin
				q			<=			16'h0000;
		end
		32'h000102C2: begin
				q			<=			16'h0000;
		end
		32'h000102C4: begin
				q			<=			16'h0000;
		end
		32'h000102C6: begin
				q			<=			16'h0000;
		end
		32'h000102C8: begin
				q			<=			16'h0000;
		end
		32'h000102CA: begin
				q			<=			16'h0000;
		end
		32'h000102CC: begin
				q			<=			16'h0000;
		end
		32'h000102CE: begin
				q			<=			16'h0000;
		end
		32'h000102D0: begin
				q			<=			16'h0000;
		end
		32'h000102D2: begin
				q			<=			16'h0000;
		end
		32'h000102D4: begin
				q			<=			16'h0000;
		end
		32'h000102D6: begin
				q			<=			16'h0000;
		end
		32'h000102D8: begin
				q			<=			16'h0000;
		end
		32'h000102DA: begin
				q			<=			16'h0000;
		end
		32'h000102DC: begin
				q			<=			16'h0000;
		end
		32'h000102DE: begin
				q			<=			16'h0000;
		end
		32'h000102E0: begin
				q			<=			16'h0000;
		end
		32'h000102E2: begin
				q			<=			16'h0000;
		end
		32'h000102E4: begin
				q			<=			16'h0000;
		end
		32'h000102E6: begin
				q			<=			16'h0000;
		end
		32'h000102E8: begin
				q			<=			16'h0000;
		end
		32'h000102EA: begin
				q			<=			16'h0000;
		end
		32'h000102EC: begin
				q			<=			16'h0000;
		end
		32'h000102EE: begin
				q			<=			16'h0000;
		end
		32'h000102F0: begin
				q			<=			16'h0000;
		end
		32'h000102F2: begin
				q			<=			16'h0000;
		end
		32'h000102F4: begin
				q			<=			16'h0000;
		end
		32'h000102F6: begin
				q			<=			16'h0000;
		end
		32'h000102F8: begin
				q			<=			16'h0000;
		end
		32'h000102FA: begin
				q			<=			16'h0000;
		end
		32'h000102FC: begin
				q			<=			16'h0000;
		end
		32'h000102FE: begin
				q			<=			16'h0000;
		end
		32'h00010300: begin
				q			<=			16'h0000;
		end
		32'h00010302: begin
				q			<=			16'h0000;
		end
		32'h00010304: begin
				q			<=			16'h0000;
		end
		32'h00010306: begin
				q			<=			16'h0000;
		end
		32'h00010308: begin
				q			<=			16'h0000;
		end
		32'h0001030A: begin
				q			<=			16'h0000;
		end
		32'h0001030C: begin
				q			<=			16'h0000;
		end
		32'h0001030E: begin
				q			<=			16'h0000;
		end
		32'h00010310: begin
				q			<=			16'h0000;
		end
		32'h00010312: begin
				q			<=			16'h0000;
		end
		32'h00010314: begin
				q			<=			16'h0000;
		end
		32'h00010316: begin
				q			<=			16'h0000;
		end
		32'h00010318: begin
				q			<=			16'h0000;
		end
		32'h0001031A: begin
				q			<=			16'h0000;
		end
		32'h0001031C: begin
				q			<=			16'h0000;
		end
		32'h0001031E: begin
				q			<=			16'h0000;
		end
		32'h00010320: begin
				q			<=			16'h0000;
		end
		32'h00010322: begin
				q			<=			16'h0000;
		end
		32'h00010324: begin
				q			<=			16'h0000;
		end
		32'h00010326: begin
				q			<=			16'h0000;
		end
		32'h00010328: begin
				q			<=			16'h0000;
		end
		32'h0001032A: begin
				q			<=			16'h0000;
		end
		32'h0001032C: begin
				q			<=			16'h0000;
		end
		32'h0001032E: begin
				q			<=			16'h0000;
		end
		32'h00010330: begin
				q			<=			16'h0000;
		end
		32'h00010332: begin
				q			<=			16'h0000;
		end
		32'h00010334: begin
				q			<=			16'h0000;
		end
		32'h00010336: begin
				q			<=			16'h0000;
		end
		32'h00010338: begin
				q			<=			16'h0000;
		end
		32'h0001033A: begin
				q			<=			16'h0000;
		end
		32'h0001033C: begin
				q			<=			16'h0000;
		end
		32'h0001033E: begin
				q			<=			16'h0000;
		end
		32'h00010340: begin
				q			<=			16'h0000;
		end
		32'h00010342: begin
				q			<=			16'h0000;
		end
		32'h00010344: begin
				q			<=			16'h0000;
		end
		32'h00010346: begin
				q			<=			16'h0000;
		end
		32'h00010348: begin
				q			<=			16'h0000;
		end
		32'h0001034A: begin
				q			<=			16'h0000;
		end
		32'h0001034C: begin
				q			<=			16'h0000;
		end
		32'h0001034E: begin
				q			<=			16'h0000;
		end
		32'h00010350: begin
				q			<=			16'h0000;
		end
		32'h00010352: begin
				q			<=			16'h0000;
		end
		32'h00010354: begin
				q			<=			16'h0000;
		end
		32'h00010356: begin
				q			<=			16'h0000;
		end
		32'h00010358: begin
				q			<=			16'h0000;
		end
		32'h0001035A: begin
				q			<=			16'h0000;
		end
		32'h0001035C: begin
				q			<=			16'h0000;
		end
		32'h0001035E: begin
				q			<=			16'h0000;
		end
		32'h00010360: begin
				q			<=			16'h0000;
		end
		32'h00010362: begin
				q			<=			16'h0000;
		end
		32'h00010364: begin
				q			<=			16'h0000;
		end
		32'h00010366: begin
				q			<=			16'h0000;
		end
		32'h00010368: begin
				q			<=			16'h0360;
		end
		32'h0001036A: begin
				q			<=			16'h0001;
		end
		32'h0001036C: begin
				q			<=			16'h0360;
		end
		32'h0001036E: begin
				q			<=			16'h0001;
		end
		32'h00010370: begin
				q			<=			16'h0368;
		end
		32'h00010372: begin
				q			<=			16'h0001;
		end
		32'h00010374: begin
				q			<=			16'h0368;
		end
		32'h00010376: begin
				q			<=			16'h0001;
		end
		32'h00010378: begin
				q			<=			16'h0370;
		end
		32'h0001037A: begin
				q			<=			16'h0001;
		end
		32'h0001037C: begin
				q			<=			16'h0370;
		end
		32'h0001037E: begin
				q			<=			16'h0001;
		end
		32'h00010380: begin
				q			<=			16'h0378;
		end
		32'h00010382: begin
				q			<=			16'h0001;
		end
		32'h00010384: begin
				q			<=			16'h0378;
		end
		32'h00010386: begin
				q			<=			16'h0001;
		end
		32'h00010388: begin
				q			<=			16'h0380;
		end
		32'h0001038A: begin
				q			<=			16'h0001;
		end
		32'h0001038C: begin
				q			<=			16'h0380;
		end
		32'h0001038E: begin
				q			<=			16'h0001;
		end
		32'h00010390: begin
				q			<=			16'h0388;
		end
		32'h00010392: begin
				q			<=			16'h0001;
		end
		32'h00010394: begin
				q			<=			16'h0388;
		end
		32'h00010396: begin
				q			<=			16'h0001;
		end
		32'h00010398: begin
				q			<=			16'h0390;
		end
		32'h0001039A: begin
				q			<=			16'h0001;
		end
		32'h0001039C: begin
				q			<=			16'h0390;
		end
		32'h0001039E: begin
				q			<=			16'h0001;
		end
		32'h000103A0: begin
				q			<=			16'h0398;
		end
		32'h000103A2: begin
				q			<=			16'h0001;
		end
		32'h000103A4: begin
				q			<=			16'h0398;
		end
		32'h000103A6: begin
				q			<=			16'h0001;
		end
		32'h000103A8: begin
				q			<=			16'h03A0;
		end
		32'h000103AA: begin
				q			<=			16'h0001;
		end
		32'h000103AC: begin
				q			<=			16'h03A0;
		end
		32'h000103AE: begin
				q			<=			16'h0001;
		end
		32'h000103B0: begin
				q			<=			16'h03A8;
		end
		32'h000103B2: begin
				q			<=			16'h0001;
		end
		32'h000103B4: begin
				q			<=			16'h03A8;
		end
		32'h000103B6: begin
				q			<=			16'h0001;
		end
		32'h000103B8: begin
				q			<=			16'h03B0;
		end
		32'h000103BA: begin
				q			<=			16'h0001;
		end
		32'h000103BC: begin
				q			<=			16'h03B0;
		end
		32'h000103BE: begin
				q			<=			16'h0001;
		end
		32'h000103C0: begin
				q			<=			16'h03B8;
		end
		32'h000103C2: begin
				q			<=			16'h0001;
		end
		32'h000103C4: begin
				q			<=			16'h03B8;
		end
		32'h000103C6: begin
				q			<=			16'h0001;
		end
		32'h000103C8: begin
				q			<=			16'h03C0;
		end
		32'h000103CA: begin
				q			<=			16'h0001;
		end
		32'h000103CC: begin
				q			<=			16'h03C0;
		end
		32'h000103CE: begin
				q			<=			16'h0001;
		end
		32'h000103D0: begin
				q			<=			16'h03C8;
		end
		32'h000103D2: begin
				q			<=			16'h0001;
		end
		32'h000103D4: begin
				q			<=			16'h03C8;
		end
		32'h000103D6: begin
				q			<=			16'h0001;
		end
		32'h000103D8: begin
				q			<=			16'h03D0;
		end
		32'h000103DA: begin
				q			<=			16'h0001;
		end
		32'h000103DC: begin
				q			<=			16'h03D0;
		end
		32'h000103DE: begin
				q			<=			16'h0001;
		end
		32'h000103E0: begin
				q			<=			16'h03D8;
		end
		32'h000103E2: begin
				q			<=			16'h0001;
		end
		32'h000103E4: begin
				q			<=			16'h03D8;
		end
		32'h000103E6: begin
				q			<=			16'h0001;
		end
		32'h000103E8: begin
				q			<=			16'h03E0;
		end
		32'h000103EA: begin
				q			<=			16'h0001;
		end
		32'h000103EC: begin
				q			<=			16'h03E0;
		end
		32'h000103EE: begin
				q			<=			16'h0001;
		end
		32'h000103F0: begin
				q			<=			16'h03E8;
		end
		32'h000103F2: begin
				q			<=			16'h0001;
		end
		32'h000103F4: begin
				q			<=			16'h03E8;
		end
		32'h000103F6: begin
				q			<=			16'h0001;
		end
		32'h000103F8: begin
				q			<=			16'h03F0;
		end
		32'h000103FA: begin
				q			<=			16'h0001;
		end
		32'h000103FC: begin
				q			<=			16'h03F0;
		end
		32'h000103FE: begin
				q			<=			16'h0001;
		end
		32'h00010400: begin
				q			<=			16'h03F8;
		end
		32'h00010402: begin
				q			<=			16'h0001;
		end
		32'h00010404: begin
				q			<=			16'h03F8;
		end
		32'h00010406: begin
				q			<=			16'h0001;
		end
		32'h00010408: begin
				q			<=			16'h0400;
		end
		32'h0001040A: begin
				q			<=			16'h0001;
		end
		32'h0001040C: begin
				q			<=			16'h0400;
		end
		32'h0001040E: begin
				q			<=			16'h0001;
		end
		32'h00010410: begin
				q			<=			16'h0408;
		end
		32'h00010412: begin
				q			<=			16'h0001;
		end
		32'h00010414: begin
				q			<=			16'h0408;
		end
		32'h00010416: begin
				q			<=			16'h0001;
		end
		32'h00010418: begin
				q			<=			16'h0410;
		end
		32'h0001041A: begin
				q			<=			16'h0001;
		end
		32'h0001041C: begin
				q			<=			16'h0410;
		end
		32'h0001041E: begin
				q			<=			16'h0001;
		end
		32'h00010420: begin
				q			<=			16'h0418;
		end
		32'h00010422: begin
				q			<=			16'h0001;
		end
		32'h00010424: begin
				q			<=			16'h0418;
		end
		32'h00010426: begin
				q			<=			16'h0001;
		end
		32'h00010428: begin
				q			<=			16'h0420;
		end
		32'h0001042A: begin
				q			<=			16'h0001;
		end
		32'h0001042C: begin
				q			<=			16'h0420;
		end
		32'h0001042E: begin
				q			<=			16'h0001;
		end
		32'h00010430: begin
				q			<=			16'h0428;
		end
		32'h00010432: begin
				q			<=			16'h0001;
		end
		32'h00010434: begin
				q			<=			16'h0428;
		end
		32'h00010436: begin
				q			<=			16'h0001;
		end
		32'h00010438: begin
				q			<=			16'h0430;
		end
		32'h0001043A: begin
				q			<=			16'h0001;
		end
		32'h0001043C: begin
				q			<=			16'h0430;
		end
		32'h0001043E: begin
				q			<=			16'h0001;
		end
		32'h00010440: begin
				q			<=			16'h0438;
		end
		32'h00010442: begin
				q			<=			16'h0001;
		end
		32'h00010444: begin
				q			<=			16'h0438;
		end
		32'h00010446: begin
				q			<=			16'h0001;
		end
		32'h00010448: begin
				q			<=			16'h0440;
		end
		32'h0001044A: begin
				q			<=			16'h0001;
		end
		32'h0001044C: begin
				q			<=			16'h0440;
		end
		32'h0001044E: begin
				q			<=			16'h0001;
		end
		32'h00010450: begin
				q			<=			16'h0448;
		end
		32'h00010452: begin
				q			<=			16'h0001;
		end
		32'h00010454: begin
				q			<=			16'h0448;
		end
		32'h00010456: begin
				q			<=			16'h0001;
		end
		32'h00010458: begin
				q			<=			16'h0450;
		end
		32'h0001045A: begin
				q			<=			16'h0001;
		end
		32'h0001045C: begin
				q			<=			16'h0450;
		end
		32'h0001045E: begin
				q			<=			16'h0001;
		end
		32'h00010460: begin
				q			<=			16'h0458;
		end
		32'h00010462: begin
				q			<=			16'h0001;
		end
		32'h00010464: begin
				q			<=			16'h0458;
		end
		32'h00010466: begin
				q			<=			16'h0001;
		end
		32'h00010468: begin
				q			<=			16'h0460;
		end
		32'h0001046A: begin
				q			<=			16'h0001;
		end
		32'h0001046C: begin
				q			<=			16'h0460;
		end
		32'h0001046E: begin
				q			<=			16'h0001;
		end
		32'h00010470: begin
				q			<=			16'h0468;
		end
		32'h00010472: begin
				q			<=			16'h0001;
		end
		32'h00010474: begin
				q			<=			16'h0468;
		end
		32'h00010476: begin
				q			<=			16'h0001;
		end
		32'h00010478: begin
				q			<=			16'h0470;
		end
		32'h0001047A: begin
				q			<=			16'h0001;
		end
		32'h0001047C: begin
				q			<=			16'h0470;
		end
		32'h0001047E: begin
				q			<=			16'h0001;
		end
		32'h00010480: begin
				q			<=			16'h0478;
		end
		32'h00010482: begin
				q			<=			16'h0001;
		end
		32'h00010484: begin
				q			<=			16'h0478;
		end
		32'h00010486: begin
				q			<=			16'h0001;
		end
		32'h00010488: begin
				q			<=			16'h0480;
		end
		32'h0001048A: begin
				q			<=			16'h0001;
		end
		32'h0001048C: begin
				q			<=			16'h0480;
		end
		32'h0001048E: begin
				q			<=			16'h0001;
		end
		32'h00010490: begin
				q			<=			16'h0488;
		end
		32'h00010492: begin
				q			<=			16'h0001;
		end
		32'h00010494: begin
				q			<=			16'h0488;
		end
		32'h00010496: begin
				q			<=			16'h0001;
		end
		32'h00010498: begin
				q			<=			16'h0490;
		end
		32'h0001049A: begin
				q			<=			16'h0001;
		end
		32'h0001049C: begin
				q			<=			16'h0490;
		end
		32'h0001049E: begin
				q			<=			16'h0001;
		end
		32'h000104A0: begin
				q			<=			16'h0498;
		end
		32'h000104A2: begin
				q			<=			16'h0001;
		end
		32'h000104A4: begin
				q			<=			16'h0498;
		end
		32'h000104A6: begin
				q			<=			16'h0001;
		end
		32'h000104A8: begin
				q			<=			16'h04A0;
		end
		32'h000104AA: begin
				q			<=			16'h0001;
		end
		32'h000104AC: begin
				q			<=			16'h04A0;
		end
		32'h000104AE: begin
				q			<=			16'h0001;
		end
		32'h000104B0: begin
				q			<=			16'h04A8;
		end
		32'h000104B2: begin
				q			<=			16'h0001;
		end
		32'h000104B4: begin
				q			<=			16'h04A8;
		end
		32'h000104B6: begin
				q			<=			16'h0001;
		end
		32'h000104B8: begin
				q			<=			16'h04B0;
		end
		32'h000104BA: begin
				q			<=			16'h0001;
		end
		32'h000104BC: begin
				q			<=			16'h04B0;
		end
		32'h000104BE: begin
				q			<=			16'h0001;
		end
		32'h000104C0: begin
				q			<=			16'h04B8;
		end
		32'h000104C2: begin
				q			<=			16'h0001;
		end
		32'h000104C4: begin
				q			<=			16'h04B8;
		end
		32'h000104C6: begin
				q			<=			16'h0001;
		end
		32'h000104C8: begin
				q			<=			16'h04C0;
		end
		32'h000104CA: begin
				q			<=			16'h0001;
		end
		32'h000104CC: begin
				q			<=			16'h04C0;
		end
		32'h000104CE: begin
				q			<=			16'h0001;
		end
		32'h000104D0: begin
				q			<=			16'h04C8;
		end
		32'h000104D2: begin
				q			<=			16'h0001;
		end
		32'h000104D4: begin
				q			<=			16'h04C8;
		end
		32'h000104D6: begin
				q			<=			16'h0001;
		end
		32'h000104D8: begin
				q			<=			16'h04D0;
		end
		32'h000104DA: begin
				q			<=			16'h0001;
		end
		32'h000104DC: begin
				q			<=			16'h04D0;
		end
		32'h000104DE: begin
				q			<=			16'h0001;
		end
		32'h000104E0: begin
				q			<=			16'h04D8;
		end
		32'h000104E2: begin
				q			<=			16'h0001;
		end
		32'h000104E4: begin
				q			<=			16'h04D8;
		end
		32'h000104E6: begin
				q			<=			16'h0001;
		end
		32'h000104E8: begin
				q			<=			16'h04E0;
		end
		32'h000104EA: begin
				q			<=			16'h0001;
		end
		32'h000104EC: begin
				q			<=			16'h04E0;
		end
		32'h000104EE: begin
				q			<=			16'h0001;
		end
		32'h000104F0: begin
				q			<=			16'h04E8;
		end
		32'h000104F2: begin
				q			<=			16'h0001;
		end
		32'h000104F4: begin
				q			<=			16'h04E8;
		end
		32'h000104F6: begin
				q			<=			16'h0001;
		end
		32'h000104F8: begin
				q			<=			16'h04F0;
		end
		32'h000104FA: begin
				q			<=			16'h0001;
		end
		32'h000104FC: begin
				q			<=			16'h04F0;
		end
		32'h000104FE: begin
				q			<=			16'h0001;
		end
		32'h00010500: begin
				q			<=			16'h04F8;
		end
		32'h00010502: begin
				q			<=			16'h0001;
		end
		32'h00010504: begin
				q			<=			16'h04F8;
		end
		32'h00010506: begin
				q			<=			16'h0001;
		end
		32'h00010508: begin
				q			<=			16'h0500;
		end
		32'h0001050A: begin
				q			<=			16'h0001;
		end
		32'h0001050C: begin
				q			<=			16'h0500;
		end
		32'h0001050E: begin
				q			<=			16'h0001;
		end
		32'h00010510: begin
				q			<=			16'h0508;
		end
		32'h00010512: begin
				q			<=			16'h0001;
		end
		32'h00010514: begin
				q			<=			16'h0508;
		end
		32'h00010516: begin
				q			<=			16'h0001;
		end
		32'h00010518: begin
				q			<=			16'h0510;
		end
		32'h0001051A: begin
				q			<=			16'h0001;
		end
		32'h0001051C: begin
				q			<=			16'h0510;
		end
		32'h0001051E: begin
				q			<=			16'h0001;
		end
		32'h00010520: begin
				q			<=			16'h0518;
		end
		32'h00010522: begin
				q			<=			16'h0001;
		end
		32'h00010524: begin
				q			<=			16'h0518;
		end
		32'h00010526: begin
				q			<=			16'h0001;
		end
		32'h00010528: begin
				q			<=			16'h0520;
		end
		32'h0001052A: begin
				q			<=			16'h0001;
		end
		32'h0001052C: begin
				q			<=			16'h0520;
		end
		32'h0001052E: begin
				q			<=			16'h0001;
		end
		32'h00010530: begin
				q			<=			16'h0528;
		end
		32'h00010532: begin
				q			<=			16'h0001;
		end
		32'h00010534: begin
				q			<=			16'h0528;
		end
		32'h00010536: begin
				q			<=			16'h0001;
		end
		32'h00010538: begin
				q			<=			16'h0530;
		end
		32'h0001053A: begin
				q			<=			16'h0001;
		end
		32'h0001053C: begin
				q			<=			16'h0530;
		end
		32'h0001053E: begin
				q			<=			16'h0001;
		end
		32'h00010540: begin
				q			<=			16'h0538;
		end
		32'h00010542: begin
				q			<=			16'h0001;
		end
		32'h00010544: begin
				q			<=			16'h0538;
		end
		32'h00010546: begin
				q			<=			16'h0001;
		end
		32'h00010548: begin
				q			<=			16'h0540;
		end
		32'h0001054A: begin
				q			<=			16'h0001;
		end
		32'h0001054C: begin
				q			<=			16'h0540;
		end
		32'h0001054E: begin
				q			<=			16'h0001;
		end
		32'h00010550: begin
				q			<=			16'h0548;
		end
		32'h00010552: begin
				q			<=			16'h0001;
		end
		32'h00010554: begin
				q			<=			16'h0548;
		end
		32'h00010556: begin
				q			<=			16'h0001;
		end
		32'h00010558: begin
				q			<=			16'h0550;
		end
		32'h0001055A: begin
				q			<=			16'h0001;
		end
		32'h0001055C: begin
				q			<=			16'h0550;
		end
		32'h0001055E: begin
				q			<=			16'h0001;
		end
		32'h00010560: begin
				q			<=			16'h0558;
		end
		32'h00010562: begin
				q			<=			16'h0001;
		end
		32'h00010564: begin
				q			<=			16'h0558;
		end
		32'h00010566: begin
				q			<=			16'h0001;
		end
		32'h00010568: begin
				q			<=			16'h0560;
		end
		32'h0001056A: begin
				q			<=			16'h0001;
		end
		32'h0001056C: begin
				q			<=			16'h0560;
		end
		32'h0001056E: begin
				q			<=			16'h0001;
		end
		32'h00010570: begin
				q			<=			16'h0568;
		end
		32'h00010572: begin
				q			<=			16'h0001;
		end
		32'h00010574: begin
				q			<=			16'h0568;
		end
		32'h00010576: begin
				q			<=			16'h0001;
		end
		32'h00010578: begin
				q			<=			16'h0570;
		end
		32'h0001057A: begin
				q			<=			16'h0001;
		end
		32'h0001057C: begin
				q			<=			16'h0570;
		end
		32'h0001057E: begin
				q			<=			16'h0001;
		end
		32'h00010580: begin
				q			<=			16'h0578;
		end
		32'h00010582: begin
				q			<=			16'h0001;
		end
		32'h00010584: begin
				q			<=			16'h0578;
		end
		32'h00010586: begin
				q			<=			16'h0001;
		end
		32'h00010588: begin
				q			<=			16'h0580;
		end
		32'h0001058A: begin
				q			<=			16'h0001;
		end
		32'h0001058C: begin
				q			<=			16'h0580;
		end
		32'h0001058E: begin
				q			<=			16'h0001;
		end
		32'h00010590: begin
				q			<=			16'h0588;
		end
		32'h00010592: begin
				q			<=			16'h0001;
		end
		32'h00010594: begin
				q			<=			16'h0588;
		end
		32'h00010596: begin
				q			<=			16'h0001;
		end
		32'h00010598: begin
				q			<=			16'h0590;
		end
		32'h0001059A: begin
				q			<=			16'h0001;
		end
		32'h0001059C: begin
				q			<=			16'h0590;
		end
		32'h0001059E: begin
				q			<=			16'h0001;
		end
		32'h000105A0: begin
				q			<=			16'h0598;
		end
		32'h000105A2: begin
				q			<=			16'h0001;
		end
		32'h000105A4: begin
				q			<=			16'h0598;
		end
		32'h000105A6: begin
				q			<=			16'h0001;
		end
		32'h000105A8: begin
				q			<=			16'h05A0;
		end
		32'h000105AA: begin
				q			<=			16'h0001;
		end
		32'h000105AC: begin
				q			<=			16'h05A0;
		end
		32'h000105AE: begin
				q			<=			16'h0001;
		end
		32'h000105B0: begin
				q			<=			16'h05A8;
		end
		32'h000105B2: begin
				q			<=			16'h0001;
		end
		32'h000105B4: begin
				q			<=			16'h05A8;
		end
		32'h000105B6: begin
				q			<=			16'h0001;
		end
		32'h000105B8: begin
				q			<=			16'h05B0;
		end
		32'h000105BA: begin
				q			<=			16'h0001;
		end
		32'h000105BC: begin
				q			<=			16'h05B0;
		end
		32'h000105BE: begin
				q			<=			16'h0001;
		end
		32'h000105C0: begin
				q			<=			16'h05B8;
		end
		32'h000105C2: begin
				q			<=			16'h0001;
		end
		32'h000105C4: begin
				q			<=			16'h05B8;
		end
		32'h000105C6: begin
				q			<=			16'h0001;
		end
		32'h000105C8: begin
				q			<=			16'h05C0;
		end
		32'h000105CA: begin
				q			<=			16'h0001;
		end
		32'h000105CC: begin
				q			<=			16'h05C0;
		end
		32'h000105CE: begin
				q			<=			16'h0001;
		end
		32'h000105D0: begin
				q			<=			16'h05C8;
		end
		32'h000105D2: begin
				q			<=			16'h0001;
		end
		32'h000105D4: begin
				q			<=			16'h05C8;
		end
		32'h000105D6: begin
				q			<=			16'h0001;
		end
		32'h000105D8: begin
				q			<=			16'h05D0;
		end
		32'h000105DA: begin
				q			<=			16'h0001;
		end
		32'h000105DC: begin
				q			<=			16'h05D0;
		end
		32'h000105DE: begin
				q			<=			16'h0001;
		end
		32'h000105E0: begin
				q			<=			16'h05D8;
		end
		32'h000105E2: begin
				q			<=			16'h0001;
		end
		32'h000105E4: begin
				q			<=			16'h05D8;
		end
		32'h000105E6: begin
				q			<=			16'h0001;
		end
		32'h000105E8: begin
				q			<=			16'h05E0;
		end
		32'h000105EA: begin
				q			<=			16'h0001;
		end
		32'h000105EC: begin
				q			<=			16'h05E0;
		end
		32'h000105EE: begin
				q			<=			16'h0001;
		end
		32'h000105F0: begin
				q			<=			16'h05E8;
		end
		32'h000105F2: begin
				q			<=			16'h0001;
		end
		32'h000105F4: begin
				q			<=			16'h05E8;
		end
		32'h000105F6: begin
				q			<=			16'h0001;
		end
		32'h000105F8: begin
				q			<=			16'h05F0;
		end
		32'h000105FA: begin
				q			<=			16'h0001;
		end
		32'h000105FC: begin
				q			<=			16'h05F0;
		end
		32'h000105FE: begin
				q			<=			16'h0001;
		end
		32'h00010600: begin
				q			<=			16'h05F8;
		end
		32'h00010602: begin
				q			<=			16'h0001;
		end
		32'h00010604: begin
				q			<=			16'h05F8;
		end
		32'h00010606: begin
				q			<=			16'h0001;
		end
		32'h00010608: begin
				q			<=			16'h0600;
		end
		32'h0001060A: begin
				q			<=			16'h0001;
		end
		32'h0001060C: begin
				q			<=			16'h0600;
		end
		32'h0001060E: begin
				q			<=			16'h0001;
		end
		32'h00010610: begin
				q			<=			16'h0608;
		end
		32'h00010612: begin
				q			<=			16'h0001;
		end
		32'h00010614: begin
				q			<=			16'h0608;
		end
		32'h00010616: begin
				q			<=			16'h0001;
		end
		32'h00010618: begin
				q			<=			16'h0610;
		end
		32'h0001061A: begin
				q			<=			16'h0001;
		end
		32'h0001061C: begin
				q			<=			16'h0610;
		end
		32'h0001061E: begin
				q			<=			16'h0001;
		end
		32'h00010620: begin
				q			<=			16'h0618;
		end
		32'h00010622: begin
				q			<=			16'h0001;
		end
		32'h00010624: begin
				q			<=			16'h0618;
		end
		32'h00010626: begin
				q			<=			16'h0001;
		end
		32'h00010628: begin
				q			<=			16'h0620;
		end
		32'h0001062A: begin
				q			<=			16'h0001;
		end
		32'h0001062C: begin
				q			<=			16'h0620;
		end
		32'h0001062E: begin
				q			<=			16'h0001;
		end
		32'h00010630: begin
				q			<=			16'h0628;
		end
		32'h00010632: begin
				q			<=			16'h0001;
		end
		32'h00010634: begin
				q			<=			16'h0628;
		end
		32'h00010636: begin
				q			<=			16'h0001;
		end
		32'h00010638: begin
				q			<=			16'h0630;
		end
		32'h0001063A: begin
				q			<=			16'h0001;
		end
		32'h0001063C: begin
				q			<=			16'h0630;
		end
		32'h0001063E: begin
				q			<=			16'h0001;
		end
		32'h00010640: begin
				q			<=			16'h0638;
		end
		32'h00010642: begin
				q			<=			16'h0001;
		end
		32'h00010644: begin
				q			<=			16'h0638;
		end
		32'h00010646: begin
				q			<=			16'h0001;
		end
		32'h00010648: begin
				q			<=			16'h0640;
		end
		32'h0001064A: begin
				q			<=			16'h0001;
		end
		32'h0001064C: begin
				q			<=			16'h0640;
		end
		32'h0001064E: begin
				q			<=			16'h0001;
		end
		32'h00010650: begin
				q			<=			16'h0648;
		end
		32'h00010652: begin
				q			<=			16'h0001;
		end
		32'h00010654: begin
				q			<=			16'h0648;
		end
		32'h00010656: begin
				q			<=			16'h0001;
		end
		32'h00010658: begin
				q			<=			16'h0650;
		end
		32'h0001065A: begin
				q			<=			16'h0001;
		end
		32'h0001065C: begin
				q			<=			16'h0650;
		end
		32'h0001065E: begin
				q			<=			16'h0001;
		end
		32'h00010660: begin
				q			<=			16'h0658;
		end
		32'h00010662: begin
				q			<=			16'h0001;
		end
		32'h00010664: begin
				q			<=			16'h0658;
		end
		32'h00010666: begin
				q			<=			16'h0001;
		end
		32'h00010668: begin
				q			<=			16'h0660;
		end
		32'h0001066A: begin
				q			<=			16'h0001;
		end
		32'h0001066C: begin
				q			<=			16'h0660;
		end
		32'h0001066E: begin
				q			<=			16'h0001;
		end
		32'h00010670: begin
				q			<=			16'h0668;
		end
		32'h00010672: begin
				q			<=			16'h0001;
		end
		32'h00010674: begin
				q			<=			16'h0668;
		end
		32'h00010676: begin
				q			<=			16'h0001;
		end
		32'h00010678: begin
				q			<=			16'h0670;
		end
		32'h0001067A: begin
				q			<=			16'h0001;
		end
		32'h0001067C: begin
				q			<=			16'h0670;
		end
		32'h0001067E: begin
				q			<=			16'h0001;
		end
		32'h00010680: begin
				q			<=			16'h0678;
		end
		32'h00010682: begin
				q			<=			16'h0001;
		end
		32'h00010684: begin
				q			<=			16'h0678;
		end
		32'h00010686: begin
				q			<=			16'h0001;
		end
		32'h00010688: begin
				q			<=			16'h0680;
		end
		32'h0001068A: begin
				q			<=			16'h0001;
		end
		32'h0001068C: begin
				q			<=			16'h0680;
		end
		32'h0001068E: begin
				q			<=			16'h0001;
		end
		32'h00010690: begin
				q			<=			16'h0688;
		end
		32'h00010692: begin
				q			<=			16'h0001;
		end
		32'h00010694: begin
				q			<=			16'h0688;
		end
		32'h00010696: begin
				q			<=			16'h0001;
		end
		32'h00010698: begin
				q			<=			16'h0690;
		end
		32'h0001069A: begin
				q			<=			16'h0001;
		end
		32'h0001069C: begin
				q			<=			16'h0690;
		end
		32'h0001069E: begin
				q			<=			16'h0001;
		end
		32'h000106A0: begin
				q			<=			16'h0698;
		end
		32'h000106A2: begin
				q			<=			16'h0001;
		end
		32'h000106A4: begin
				q			<=			16'h0698;
		end
		32'h000106A6: begin
				q			<=			16'h0001;
		end
		32'h000106A8: begin
				q			<=			16'h06A0;
		end
		32'h000106AA: begin
				q			<=			16'h0001;
		end
		32'h000106AC: begin
				q			<=			16'h06A0;
		end
		32'h000106AE: begin
				q			<=			16'h0001;
		end
		32'h000106B0: begin
				q			<=			16'h06A8;
		end
		32'h000106B2: begin
				q			<=			16'h0001;
		end
		32'h000106B4: begin
				q			<=			16'h06A8;
		end
		32'h000106B6: begin
				q			<=			16'h0001;
		end
		32'h000106B8: begin
				q			<=			16'h06B0;
		end
		32'h000106BA: begin
				q			<=			16'h0001;
		end
		32'h000106BC: begin
				q			<=			16'h06B0;
		end
		32'h000106BE: begin
				q			<=			16'h0001;
		end
		32'h000106C0: begin
				q			<=			16'h06B8;
		end
		32'h000106C2: begin
				q			<=			16'h0001;
		end
		32'h000106C4: begin
				q			<=			16'h06B8;
		end
		32'h000106C6: begin
				q			<=			16'h0001;
		end
		32'h000106C8: begin
				q			<=			16'h06C0;
		end
		32'h000106CA: begin
				q			<=			16'h0001;
		end
		32'h000106CC: begin
				q			<=			16'h06C0;
		end
		32'h000106CE: begin
				q			<=			16'h0001;
		end
		32'h000106D0: begin
				q			<=			16'h06C8;
		end
		32'h000106D2: begin
				q			<=			16'h0001;
		end
		32'h000106D4: begin
				q			<=			16'h06C8;
		end
		32'h000106D6: begin
				q			<=			16'h0001;
		end
		32'h000106D8: begin
				q			<=			16'h06D0;
		end
		32'h000106DA: begin
				q			<=			16'h0001;
		end
		32'h000106DC: begin
				q			<=			16'h06D0;
		end
		32'h000106DE: begin
				q			<=			16'h0001;
		end
		32'h000106E0: begin
				q			<=			16'h06D8;
		end
		32'h000106E2: begin
				q			<=			16'h0001;
		end
		32'h000106E4: begin
				q			<=			16'h06D8;
		end
		32'h000106E6: begin
				q			<=			16'h0001;
		end
		32'h000106E8: begin
				q			<=			16'h06E0;
		end
		32'h000106EA: begin
				q			<=			16'h0001;
		end
		32'h000106EC: begin
				q			<=			16'h06E0;
		end
		32'h000106EE: begin
				q			<=			16'h0001;
		end
		32'h000106F0: begin
				q			<=			16'h06E8;
		end
		32'h000106F2: begin
				q			<=			16'h0001;
		end
		32'h000106F4: begin
				q			<=			16'h06E8;
		end
		32'h000106F6: begin
				q			<=			16'h0001;
		end
		32'h000106F8: begin
				q			<=			16'h06F0;
		end
		32'h000106FA: begin
				q			<=			16'h0001;
		end
		32'h000106FC: begin
				q			<=			16'h06F0;
		end
		32'h000106FE: begin
				q			<=			16'h0001;
		end
		32'h00010700: begin
				q			<=			16'h06F8;
		end
		32'h00010702: begin
				q			<=			16'h0001;
		end
		32'h00010704: begin
				q			<=			16'h06F8;
		end
		32'h00010706: begin
				q			<=			16'h0001;
		end
		32'h00010708: begin
				q			<=			16'h0700;
		end
		32'h0001070A: begin
				q			<=			16'h0001;
		end
		32'h0001070C: begin
				q			<=			16'h0700;
		end
		32'h0001070E: begin
				q			<=			16'h0001;
		end
		32'h00010710: begin
				q			<=			16'h0708;
		end
		32'h00010712: begin
				q			<=			16'h0001;
		end
		32'h00010714: begin
				q			<=			16'h0708;
		end
		32'h00010716: begin
				q			<=			16'h0001;
		end
		32'h00010718: begin
				q			<=			16'h0710;
		end
		32'h0001071A: begin
				q			<=			16'h0001;
		end
		32'h0001071C: begin
				q			<=			16'h0710;
		end
		32'h0001071E: begin
				q			<=			16'h0001;
		end
		32'h00010720: begin
				q			<=			16'h0718;
		end
		32'h00010722: begin
				q			<=			16'h0001;
		end
		32'h00010724: begin
				q			<=			16'h0718;
		end
		32'h00010726: begin
				q			<=			16'h0001;
		end
		32'h00010728: begin
				q			<=			16'h0720;
		end
		32'h0001072A: begin
				q			<=			16'h0001;
		end
		32'h0001072C: begin
				q			<=			16'h0720;
		end
		32'h0001072E: begin
				q			<=			16'h0001;
		end
		32'h00010730: begin
				q			<=			16'h0728;
		end
		32'h00010732: begin
				q			<=			16'h0001;
		end
		32'h00010734: begin
				q			<=			16'h0728;
		end
		32'h00010736: begin
				q			<=			16'h0001;
		end
		32'h00010738: begin
				q			<=			16'h0730;
		end
		32'h0001073A: begin
				q			<=			16'h0001;
		end
		32'h0001073C: begin
				q			<=			16'h0730;
		end
		32'h0001073E: begin
				q			<=			16'h0001;
		end
		32'h00010740: begin
				q			<=			16'h0738;
		end
		32'h00010742: begin
				q			<=			16'h0001;
		end
		32'h00010744: begin
				q			<=			16'h0738;
		end
		32'h00010746: begin
				q			<=			16'h0001;
		end
		32'h00010748: begin
				q			<=			16'h0740;
		end
		32'h0001074A: begin
				q			<=			16'h0001;
		end
		32'h0001074C: begin
				q			<=			16'h0740;
		end
		32'h0001074E: begin
				q			<=			16'h0001;
		end
		32'h00010750: begin
				q			<=			16'h0748;
		end
		32'h00010752: begin
				q			<=			16'h0001;
		end
		32'h00010754: begin
				q			<=			16'h0748;
		end
		32'h00010756: begin
				q			<=			16'h0001;
		end
		32'h00010758: begin
				q			<=			16'h0750;
		end
		32'h0001075A: begin
				q			<=			16'h0001;
		end
		32'h0001075C: begin
				q			<=			16'h0750;
		end
		32'h0001075E: begin
				q			<=			16'h0001;
		end
		32'h00010760: begin
				q			<=			16'h0758;
		end
		32'h00010762: begin
				q			<=			16'h0001;
		end
		32'h00010764: begin
				q			<=			16'h0758;
		end
		32'h00010766: begin
				q			<=			16'h0001;
		end
		32'h00010768: begin
				q			<=			16'h0043;
		end
		32'h0001076A: begin
				q			<=			16'h0000;
		end
		32'h0001076C: begin
				q			<=			16'h0000;
		end
		32'h0001076E: begin
				q			<=			16'h0000;
		end
		32'h00010770: begin
				q			<=			16'h0000;
		end
		32'h00010772: begin
				q			<=			16'h0000;
		end
		32'h00010774: begin
				q			<=			16'h0000;
		end
		32'h00010776: begin
				q			<=			16'h0000;
		end
		32'h00010778: begin
				q			<=			16'h0000;
		end
		32'h0001077A: begin
				q			<=			16'h0000;
		end
		32'h0001077C: begin
				q			<=			16'h0000;
		end
		32'h0001077E: begin
				q			<=			16'h0000;
		end
		32'h00010780: begin
				q			<=			16'h0000;
		end
		32'h00010782: begin
				q			<=			16'h0000;
		end
		32'h00010784: begin
				q			<=			16'h0000;
		end
		32'h00010786: begin
				q			<=			16'h0000;
		end
		32'h00010788: begin
				q			<=			16'h0043;
		end
		32'h0001078A: begin
				q			<=			16'h0000;
		end
		32'h0001078C: begin
				q			<=			16'h0000;
		end
		32'h0001078E: begin
				q			<=			16'h0000;
		end
		32'h00010790: begin
				q			<=			16'h0000;
		end
		32'h00010792: begin
				q			<=			16'h0000;
		end
		32'h00010794: begin
				q			<=			16'h0000;
		end
		32'h00010796: begin
				q			<=			16'h0000;
		end
		32'h00010798: begin
				q			<=			16'h0000;
		end
		32'h0001079A: begin
				q			<=			16'h0000;
		end
		32'h0001079C: begin
				q			<=			16'h0000;
		end
		32'h0001079E: begin
				q			<=			16'h0000;
		end
		32'h000107A0: begin
				q			<=			16'h0000;
		end
		32'h000107A2: begin
				q			<=			16'h0000;
		end
		32'h000107A4: begin
				q			<=			16'h0000;
		end
		32'h000107A6: begin
				q			<=			16'h0000;
		end
		32'h000107A8: begin
				q			<=			16'h0043;
		end
		32'h000107AA: begin
				q			<=			16'h0000;
		end
		32'h000107AC: begin
				q			<=			16'h0000;
		end
		32'h000107AE: begin
				q			<=			16'h0000;
		end
		32'h000107B0: begin
				q			<=			16'h0000;
		end
		32'h000107B2: begin
				q			<=			16'h0000;
		end
		32'h000107B4: begin
				q			<=			16'h0000;
		end
		32'h000107B6: begin
				q			<=			16'h0000;
		end
		32'h000107B8: begin
				q			<=			16'h0000;
		end
		32'h000107BA: begin
				q			<=			16'h0000;
		end
		32'h000107BC: begin
				q			<=			16'h0000;
		end
		32'h000107BE: begin
				q			<=			16'h0000;
		end
		32'h000107C0: begin
				q			<=			16'h0000;
		end
		32'h000107C2: begin
				q			<=			16'h0000;
		end
		32'h000107C4: begin
				q			<=			16'h0000;
		end
		32'h000107C6: begin
				q			<=			16'h0000;
		end
		32'h000107C8: begin
				q			<=			16'h0043;
		end
		32'h000107CA: begin
				q			<=			16'h0000;
		end
		32'h000107CC: begin
				q			<=			16'h0000;
		end
		32'h000107CE: begin
				q			<=			16'h0000;
		end
		32'h000107D0: begin
				q			<=			16'h0000;
		end
		32'h000107D2: begin
				q			<=			16'h0000;
		end
		32'h000107D4: begin
				q			<=			16'h0000;
		end
		32'h000107D6: begin
				q			<=			16'h0000;
		end
		32'h000107D8: begin
				q			<=			16'h0000;
		end
		32'h000107DA: begin
				q			<=			16'h0000;
		end
		32'h000107DC: begin
				q			<=			16'h0000;
		end
		32'h000107DE: begin
				q			<=			16'h0000;
		end
		32'h000107E0: begin
				q			<=			16'h0000;
		end
		32'h000107E2: begin
				q			<=			16'h0000;
		end
		32'h000107E4: begin
				q			<=			16'h0000;
		end
		32'h000107E6: begin
				q			<=			16'h0000;
		end
		32'h000107E8: begin
				q			<=			16'h0043;
		end
		32'h000107EA: begin
				q			<=			16'h0000;
		end
		32'h000107EC: begin
				q			<=			16'h0000;
		end
		32'h000107EE: begin
				q			<=			16'h0000;
		end
		32'h000107F0: begin
				q			<=			16'h0000;
		end
		32'h000107F2: begin
				q			<=			16'h0000;
		end
		32'h000107F4: begin
				q			<=			16'h0000;
		end
		32'h000107F6: begin
				q			<=			16'h0000;
		end
		32'h000107F8: begin
				q			<=			16'h0000;
		end
		32'h000107FA: begin
				q			<=			16'h0000;
		end
		32'h000107FC: begin
				q			<=			16'h0000;
		end
		32'h000107FE: begin
				q			<=			16'h0000;
		end
		32'h00010800: begin
				q			<=			16'h0000;
		end
		32'h00010802: begin
				q			<=			16'h0000;
		end
		32'h00010804: begin
				q			<=			16'h0000;
		end
		32'h00010806: begin
				q			<=			16'h0000;
		end
		32'h00010808: begin
				q			<=			16'h0043;
		end
		32'h0001080A: begin
				q			<=			16'h0000;
		end
		32'h0001080C: begin
				q			<=			16'h0000;
		end
		32'h0001080E: begin
				q			<=			16'h0000;
		end
		32'h00010810: begin
				q			<=			16'h0000;
		end
		32'h00010812: begin
				q			<=			16'h0000;
		end
		32'h00010814: begin
				q			<=			16'h0000;
		end
		32'h00010816: begin
				q			<=			16'h0000;
		end
		32'h00010818: begin
				q			<=			16'h0000;
		end
		32'h0001081A: begin
				q			<=			16'h0000;
		end
		32'h0001081C: begin
				q			<=			16'h0000;
		end
		32'h0001081E: begin
				q			<=			16'h0000;
		end
		32'h00010820: begin
				q			<=			16'h0000;
		end
		32'h00010822: begin
				q			<=			16'h0000;
		end
		32'h00010824: begin
				q			<=			16'h0000;
		end
		32'h00010826: begin
				q			<=			16'h0000;
		end
		32'h00010828: begin
				q			<=			16'h0043;
		end
		32'h0001082A: begin
				q			<=			16'h0000;
		end
		32'h0001082C: begin
				q			<=			16'h0000;
		end
		32'h0001082E: begin
				q			<=			16'h0000;
		end
		32'h00010830: begin
				q			<=			16'h0000;
		end
		32'h00010832: begin
				q			<=			16'h0000;
		end
		32'h00010834: begin
				q			<=			16'h0000;
		end
		32'h00010836: begin
				q			<=			16'h0000;
		end
		32'h00010838: begin
				q			<=			16'h0000;
		end
		32'h0001083A: begin
				q			<=			16'h0000;
		end
		32'h0001083C: begin
				q			<=			16'h0000;
		end
		32'h0001083E: begin
				q			<=			16'h0000;
		end
		32'h00010840: begin
				q			<=			16'h0000;
		end
		32'h00010842: begin
				q			<=			16'h0000;
		end
		32'h00010844: begin
				q			<=			16'h0000;
		end
		32'h00010846: begin
				q			<=			16'h0000;
		end
		32'h00010848: begin
				q			<=			16'hA49C;
		end
		32'h0001084A: begin
				q			<=			16'h0000;
		end
		32'h0001084C: begin
				q			<=			16'h9B7C;
		end
		32'h0001084E: begin
				q			<=			16'h0000;
		end
		32'h00010850: begin
				q			<=			16'h0000;
		end
		32'h00010852: begin
				q			<=			16'h0000;
		end
		32'h00010854: begin
				q			<=			16'hF7B4;
		end
		32'h00010856: begin
				q			<=			16'h0000;
		end
		32'h00010858: begin
				q			<=			16'hFDE4;
		end
		32'h0001085A: begin
				q			<=			16'h0000;
		end
		32'h0001085C: begin
				q			<=			16'hFDA8;
		end
		32'h0001085E: begin
				q			<=			16'h0000;
		end
		32'h00010860: begin
				q			<=			16'hFDA8;
		end
		32'h00010862: begin
				q			<=			16'h0000;
		end
		32'h00010864: begin
				q			<=			16'hFDA8;
		end
		32'h00010866: begin
				q			<=			16'h0000;
		end
		32'h00010868: begin
				q			<=			16'hFDA8;
		end
		32'h0001086A: begin
				q			<=			16'h0000;
		end
		32'h0001086C: begin
				q			<=			16'hFDA8;
		end
		32'h0001086E: begin
				q			<=			16'h0000;
		end
		32'h00010870: begin
				q			<=			16'hFDA8;
		end
		32'h00010872: begin
				q			<=			16'h0000;
		end
		32'h00010874: begin
				q			<=			16'hFDA8;
		end
		32'h00010876: begin
				q			<=			16'h0000;
		end
		32'h00010878: begin
				q			<=			16'hFDA8;
		end
		32'h0001087A: begin
				q			<=			16'h0000;
		end
		32'h0001087C: begin
				q			<=			16'hFDA8;
		end
		32'h0001087E: begin
				q			<=			16'h0000;
		end
		32'h00010880: begin
				q			<=			16'hFFFF;
		end
		32'h00010882: begin
				q			<=			16'hFFFF;
		end
		32'h00010884: begin
				q			<=			16'hFFFF;
		end
		32'h00010886: begin
				q			<=			16'hFFFF;
		end
		32'h00010888: begin
				q			<=			16'hFFFF;
		end
		32'h0001088A: begin
				q			<=			16'hFFFF;
		end
		32'h0001088C: begin
				q			<=			16'hFFFF;
		end
		32'h0001088E: begin
				q			<=			16'h0000;
		end
		32'h00010890: begin
				q			<=			16'h0001;
		end
		32'h00010892: begin
				q			<=			16'h5341;
		end
		32'h00010894: begin
				q			<=			16'h4943;
		end
		32'h00010896: begin
				q			<=			16'h0049;
		end
		32'h00010898: begin
				q			<=			16'h0000;
		end
		32'h0001089A: begin
				q			<=			16'h0000;
		end
		32'h0001089C: begin
				q			<=			16'h0000;
		end
		32'h0001089E: begin
				q			<=			16'h0000;
		end
		32'h000108A0: begin
				q			<=			16'h0000;
		end
		32'h000108A2: begin
				q			<=			16'h0000;
		end
		32'h000108A4: begin
				q			<=			16'h0000;
		end
		32'h000108A6: begin
				q			<=			16'h0000;
		end
		32'h000108A8: begin
				q			<=			16'h0000;
		end
		32'h000108AA: begin
				q			<=			16'h0000;
		end
		32'h000108AC: begin
				q			<=			16'h0000;
		end
		32'h000108AE: begin
				q			<=			16'h0000;
		end
		32'h000108B0: begin
				q			<=			16'h0000;
		end
		32'h000108B2: begin
				q			<=			16'h5341;
		end
		32'h000108B4: begin
				q			<=			16'h4943;
		end
		32'h000108B6: begin
				q			<=			16'h0049;
		end
		32'h000108B8: begin
				q			<=			16'h0000;
		end
		32'h000108BA: begin
				q			<=			16'h0000;
		end
		32'h000108BC: begin
				q			<=			16'h0000;
		end
		32'h000108BE: begin
				q			<=			16'h0000;
		end
		32'h000108C0: begin
				q			<=			16'h0000;
		end
		32'h000108C2: begin
				q			<=			16'h0000;
		end
		32'h000108C4: begin
				q			<=			16'h0000;
		end
		32'h000108C6: begin
				q			<=			16'h0000;
		end
		32'h000108C8: begin
				q			<=			16'h0000;
		end
		32'h000108CA: begin
				q			<=			16'h0000;
		end
		32'h000108CC: begin
				q			<=			16'h0000;
		end
		32'h000108CE: begin
				q			<=			16'h0000;
		end
		32'h000108D0: begin
				q			<=			16'h0000;
		end
		32'h000108D2: begin
				q			<=			16'h0000;
		end
		32'h000108D4: begin
				q			<=			16'hFF38;
		end
		32'h000108D6: begin
				q			<=			16'h0000;
		end
		32'h000108D8: begin
				q			<=			16'hFF38;
		end
		32'h000108DA: begin
				q			<=			16'h0000;
		end
		32'h000108DC: begin
				q			<=			16'hFFFF;
		end
		32'h000108DE: begin
				q			<=			16'hFFFF;
		end
		32'h000108E0: begin
				q			<=			16'h0000;
		end
		32'h000108E2: begin
				q			<=			16'h0002;
		end
		32'h000108E4: begin
				q			<=			16'h0031;
		end
		32'h000108E6: begin
				q			<=			16'h0000;
		end
		32'h000108E8: begin
				q			<=			16'h0030;
		end
		32'h000108EA: begin
				q			<=			16'h0000;
		end
		32'h000108EC: begin
				q			<=			16'h0000;
		end
		32'h000108EE: begin
				q			<=			16'h0100;
		end
		32'h000108F0: begin
				q			<=			16'hFFFF;
		end
		32'h000108F2: begin
				q			<=			16'h1FFF;
		end
		default: begin
				q			<=			16'h0000;
		end
	endcase
end

endmodule

////////////////////////////////////////////////////////
// GERANIUM SYSTEM INCLUDE										//
////////////////////////////////////////////////////////

`timescale 1ps / 1ps

`ifndef INCLUDE_SYSTEM
`define INCLUDE_SYSTEM 1

///////////////////////////////////////////////////////////////////////
// CONSTANTS																			//
///////////////////////////////////////////////////////////////////////

parameter TOTAL_DMA_CHANNELS					=		1;

///////////////////////////////////////////////////////////////////////
// DMA STRUCTS																			//
///////////////////////////////////////////////////////////////////////

typedef
struct
packed
{
	logic		[27:0]		addr;
	logic						setaddr;
	logic		[31:0]		reqlen;
	logic						setreqlen;
	logic						req;
	logic						active;

} dma_channel_fromhost;

typedef
struct
packed
{
	logic						valid;
	logic		[15:0]		data;
	
} dma_channel_tohost;

///////////////////////////////////////////////////////////////////////
// TYPEDEFS																				//
///////////////////////////////////////////////////////////////////////

typedef dma_channel_fromhost				[TOTAL_DMA_CHANNELS-1:0]														dma_channels_from_host;
typedef dma_channel_tohost					[TOTAL_DMA_CHANNELS-1:0]														dma_channels_to_host;

`endif
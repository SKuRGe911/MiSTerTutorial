// avalonslavetestbench.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module avalonslavetestbench (
		input  wire [63:0] avalon_writedata,     // avalon.writedata
		input  wire [7:0]  avalon_burstcount,    //       .burstcount
		output wire [63:0] avalon_readdata,      //       .readdata
		input  wire [28:0] avalon_address,       //       .address
		output wire        avalon_waitrequest,   //       .waitrequest
		input  wire        avalon_write,         //       .write
		input  wire        avalon_read,          //       .read
		input  wire [7:0]  avalon_byteenable,    //       .byteenable
		output wire        avalon_readdatavalid, //       .readdatavalid
		input  wire        clk_clk,              //    clk.clk
		input  wire        reset_reset           //  reset.reset
	);

	altera_avalon_mm_slave_bfm #(
		.AV_ADDRESS_W               (29),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (8),
		.AV_BURSTCOUNT_W            (8),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (1),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) mm_slave_bfm_0 (
		.clk                      (clk_clk),              //       clk.clk
		.reset                    (reset_reset),          // clk_reset.reset
		.avs_writedata            (avalon_writedata),     //        s0.writedata
		.avs_burstcount           (avalon_burstcount),    //          .burstcount
		.avs_readdata             (avalon_readdata),      //          .readdata
		.avs_address              (avalon_address),       //          .address
		.avs_waitrequest          (avalon_waitrequest),   //          .waitrequest
		.avs_write                (avalon_write),         //          .write
		.avs_read                 (avalon_read),          //          .read
		.avs_byteenable           (avalon_byteenable),    //          .byteenable
		.avs_readdatavalid        (avalon_readdatavalid), //          .readdatavalid
		.avs_begintransfer        (1'b0),                 // (terminated)
		.avs_beginbursttransfer   (1'b0),                 // (terminated)
		.avs_arbiterlock          (1'b0),                 // (terminated)
		.avs_lock                 (1'b0),                 // (terminated)
		.avs_debugaccess          (1'b0),                 // (terminated)
		.avs_transactionid        (8'b00000000),          // (terminated)
		.avs_readid               (),                     // (terminated)
		.avs_writeid              (),                     // (terminated)
		.avs_clken                (1'b1),                 // (terminated)
		.avs_response             (),                     // (terminated)
		.avs_writeresponserequest (1'b0),                 // (terminated)
		.avs_writeresponsevalid   (),                     // (terminated)
		.avs_readresponse         (),                     // (terminated)
		.avs_writeresponse        ()                      // (terminated)
	);

endmodule
